--------------------------------------------------------------------------
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bramMacro is
   port(
      clka: in std_logic;        -- data
      clkb: in std_logic;        -- vga
      a_addr : in std_logic_vector(11 downto 0);
      b_addr: in std_logic_vector(11 downto 0);
      a_we : in std_logic;
      a_din : in std_logic_vector(7 downto 0);
      a_dout : out std_logic_vector(7 downto 0);
      b_dout : out std_logic_vector(7 downto 0)
   );
end bramMacro;

architecture arch of bramMacro is
    -- 64 zeros: 64 x 4 = 256
	constant INIT_VAL_256 : bit_Vector(255 downto 0) :=
    X"0000000000000000000000000000000000000000000000000000000000000000";
    constant INIT_VAL_36 : bit_Vector(255 downto 0) := X"000000000";

----- component RAMB36E1 -----
component RAMB36E1
  generic (
     DOA_REG : integer := 0;
     DOB_REG : integer := 0;
     EN_ECC_READ : boolean := FALSE;
     EN_ECC_WRITE : boolean := FALSE;
     INITP_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INITP_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_00 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_01 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_02 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_03 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_04 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_05 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_06 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_07 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_08 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_09 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_0F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_10 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_11 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_12 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_13 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_14 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_15 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_16 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_17 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_18 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_19 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_1F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_20 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_21 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_22 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_23 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_24 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_25 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_26 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_27 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_28 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_29 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_2F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_30 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_31 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_32 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_33 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_34 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_35 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_36 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_37 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_38 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_39 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_3F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_40 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_41 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_42 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_43 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_44 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_45 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_46 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_47 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_48 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_49 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_4F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_50 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_51 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_52 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_53 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_54 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_55 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_56 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_57 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_58 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_59 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_5F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_60 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_61 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_62 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_63 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_64 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_65 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_66 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_67 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_68 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_69 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_6F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_70 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_71 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_72 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_73 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_74 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_75 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_76 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_77 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_78 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_79 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_7F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
     INIT_A : bit_vector := X"000000000";
     INIT_B : bit_vector := X"000000000";
     INIT_FILE : string := "NONE";
     IS_CLKARDCLK_INVERTED : bit := '0';
     IS_CLKBWRCLK_INVERTED : bit := '0';
     IS_ENARDEN_INVERTED : bit := '0';
     IS_ENBWREN_INVERTED : bit := '0';
     IS_RSTRAMARSTRAM_INVERTED : bit := '0';
     IS_RSTRAMB_INVERTED : bit := '0';
     IS_RSTREGARSTREG_INVERTED : bit := '0';
     IS_RSTREGB_INVERTED : bit := '0';
     RAM_EXTENSION_A : string := "NONE";
     RAM_EXTENSION_B : string := "NONE";
     RAM_MODE : string := "TDP";
     RDADDR_COLLISION_HWCONFIG : string := "DELAYED_WRITE";
     READ_WIDTH_A : integer := 0;
     READ_WIDTH_B : integer := 0;
     RSTREG_PRIORITY_A : string := "RSTREG";
     RSTREG_PRIORITY_B : string := "RSTREG";
     SIM_COLLISION_CHECK : string := "ALL";
     SIM_DEVICE : string := "7SERIES";
     SRVAL_A : bit_vector := X"000000000";
     SRVAL_B : bit_vector := X"000000000";
     WRITE_MODE_A : string := "WRITE_FIRST";
     WRITE_MODE_B : string := "WRITE_FIRST";
     WRITE_WIDTH_A : integer := 0;
     WRITE_WIDTH_B : integer := 0
  );
  port (
     CASCADEOUTA : out std_ulogic;
     CASCADEOUTB : out std_ulogic;
     DBITERR : out std_ulogic;
     DOADO : out std_logic_vector(31 downto 0);
     DOBDO : out std_logic_vector(31 downto 0);
     DOPADOP : out std_logic_vector(3 downto 0);
     DOPBDOP : out std_logic_vector(3 downto 0);
     ECCPARITY : out std_logic_vector(7 downto 0);
     RDADDRECC : out std_logic_vector(8 downto 0);
     SBITERR : out std_ulogic;
     ADDRARDADDR : in std_logic_vector(15 downto 0);
     ADDRBWRADDR : in std_logic_vector(15 downto 0);
     CASCADEINA : in std_ulogic;
     CASCADEINB : in std_ulogic;
     CLKARDCLK : in std_ulogic;
     CLKBWRCLK : in std_ulogic;
     DIADI : in std_logic_vector(31 downto 0);
     DIBDI : in std_logic_vector(31 downto 0);
     DIPADIP : in std_logic_vector(3 downto 0);
     DIPBDIP : in std_logic_vector(3 downto 0);
     ENARDEN : in std_ulogic;
     ENBWREN : in std_ulogic;
     INJECTDBITERR : in std_ulogic;
     INJECTSBITERR : in std_ulogic;
     REGCEAREGCE : in std_ulogic;
     REGCEB : in std_ulogic;
     RSTRAMARSTRAM : in std_ulogic;
     RSTRAMB : in std_ulogic;
     RSTREGARSTREG : in std_ulogic;
     RSTREGB : in std_ulogic;
     WEA : in std_logic_vector(3 downto 0);
     WEBWE : in std_logic_vector(7 downto 0)
  );
end component;

begin

  BRAM_inst : RAMB36E1
  generic map (
    DOA_REG => 0,
    DOB_REG => 0,
    EN_ECC_READ => FALSE,
    EN_ECC_WRITE => FALSE,
      INITP_00 => INIT_VAL_256,
      INITP_01 => INIT_VAL_256,
      INITP_02 => INIT_VAL_256,
      INITP_03 => INIT_VAL_256,
      INITP_04 => INIT_VAL_256,
      INITP_05 => INIT_VAL_256,
      INITP_06 => INIT_VAL_256,
      INITP_07 => INIT_VAL_256,
      INITP_08 => INIT_VAL_256,
      INITP_09 => INIT_VAL_256,
      INITP_0A => INIT_VAL_256,
      INITP_0B => INIT_VAL_256,
      INITP_0C => INIT_VAL_256,
      INITP_0D => INIT_VAL_256,
      INITP_0E => INIT_VAL_256,
      INITP_0F => INIT_VAL_256,
      INIT_00 => INIT_VAL_256,
      INIT_01 => INIT_VAL_256,
      INIT_02 => INIT_VAL_256,
      INIT_03 => INIT_VAL_256,
      INIT_04 => INIT_VAL_256,
      INIT_05 => INIT_VAL_256,
      INIT_06 => INIT_VAL_256,
      INIT_07 => INIT_VAL_256,
      INIT_08 => INIT_VAL_256,
      INIT_09 => INIT_VAL_256,
      INIT_0A => INIT_VAL_256,
      INIT_0B => INIT_VAL_256,
      INIT_0C => INIT_VAL_256,
      INIT_0D => INIT_VAL_256,
      INIT_0E => INIT_VAL_256,
      INIT_0F => INIT_VAL_256,
      INIT_10 => INIT_VAL_256,
      INIT_11 => INIT_VAL_256,
      INIT_12 => INIT_VAL_256,
      INIT_13 => INIT_VAL_256,
      INIT_14 => INIT_VAL_256,
      INIT_15 => INIT_VAL_256,
      INIT_16 => INIT_VAL_256,
      INIT_17 => INIT_VAL_256,
      INIT_18 => INIT_VAL_256,
      INIT_19 => INIT_VAL_256,
      INIT_1A => INIT_VAL_256,
      INIT_1B => INIT_VAL_256,
      INIT_1C => INIT_VAL_256,
      INIT_1D => INIT_VAL_256,
      INIT_1E => INIT_VAL_256,
      INIT_1F => INIT_VAL_256,
      INIT_20 => INIT_VAL_256,
      INIT_21 => INIT_VAL_256,
      INIT_22 => INIT_VAL_256,
      INIT_23 => INIT_VAL_256,
      INIT_24 => INIT_VAL_256,
      INIT_25 => INIT_VAL_256,
      INIT_26 => INIT_VAL_256,
      INIT_27 => INIT_VAL_256,
      INIT_28 => INIT_VAL_256,
      INIT_29 => INIT_VAL_256,
      INIT_2A => INIT_VAL_256,
      INIT_2B => INIT_VAL_256,
      INIT_2C => INIT_VAL_256,
      INIT_2D => INIT_VAL_256,
      INIT_2E => INIT_VAL_256,
      INIT_2F => INIT_VAL_256,
      INIT_30 => INIT_VAL_256,
      INIT_31 => INIT_VAL_256,
      INIT_32 => INIT_VAL_256,
      INIT_33 => INIT_VAL_256,
      INIT_34 => INIT_VAL_256,
      INIT_35 => INIT_VAL_256,
      INIT_36 => INIT_VAL_256,
      INIT_37 => INIT_VAL_256,
      INIT_38 => INIT_VAL_256,
      INIT_39 => INIT_VAL_256,
      INIT_3A => INIT_VAL_256,
      INIT_3B => INIT_VAL_256,
      INIT_3C => INIT_VAL_256,
      INIT_3D => INIT_VAL_256,
      INIT_3E => INIT_VAL_256,
      INIT_3F => INIT_VAL_256,
      INIT_40 => INIT_VAL_256,
      INIT_41 => INIT_VAL_256,
      INIT_42 => INIT_VAL_256,
      INIT_43 => INIT_VAL_256,
      INIT_44 => INIT_VAL_256,
      INIT_45 => INIT_VAL_256,
      INIT_46 => INIT_VAL_256,
      INIT_47 => INIT_VAL_256,
      INIT_48 => INIT_VAL_256,
      INIT_49 => INIT_VAL_256,
      INIT_4A => INIT_VAL_256,
      INIT_4B => INIT_VAL_256,
      INIT_4C => INIT_VAL_256,
      INIT_4D => INIT_VAL_256,
      INIT_4E => INIT_VAL_256,
      INIT_4F => INIT_VAL_256,
      INIT_50 => INIT_VAL_256,
      INIT_51 => INIT_VAL_256,
      INIT_52 => INIT_VAL_256,
      INIT_53 => INIT_VAL_256,
      INIT_54 => INIT_VAL_256,
      INIT_55 => INIT_VAL_256,
      INIT_56 => INIT_VAL_256,
      INIT_57 => INIT_VAL_256,
      INIT_58 => INIT_VAL_256,
      INIT_59 => INIT_VAL_256,
      INIT_5A => INIT_VAL_256,
      INIT_5B => INIT_VAL_256,
      INIT_5C => INIT_VAL_256,
      INIT_5D => INIT_VAL_256,
      INIT_5E => INIT_VAL_256,
      INIT_5F => INIT_VAL_256,
      INIT_60 => INIT_VAL_256,
      INIT_61 => INIT_VAL_256,
      INIT_62 => INIT_VAL_256,
      INIT_63 => INIT_VAL_256,
      INIT_64 => INIT_VAL_256,
      INIT_65 => INIT_VAL_256,
      INIT_66 => INIT_VAL_256,
      INIT_67 => INIT_VAL_256,
      INIT_68 => INIT_VAL_256,
      INIT_69 => INIT_VAL_256,
      INIT_6A => INIT_VAL_256,
      INIT_6B => INIT_VAL_256,
      INIT_6C => INIT_VAL_256,
      INIT_6D => INIT_VAL_256,
      INIT_6E => INIT_VAL_256,
      INIT_6F => INIT_VAL_256,
      INIT_70 => INIT_VAL_256,
      INIT_71 => INIT_VAL_256,
      INIT_72 => INIT_VAL_256,
      INIT_73 => INIT_VAL_256,
      INIT_74 => INIT_VAL_256,
      INIT_75 => INIT_VAL_256,
      INIT_76 => INIT_VAL_256,
      INIT_77 => INIT_VAL_256,
      INIT_78 => INIT_VAL_256,
      INIT_79 => INIT_VAL_256,
      INIT_7A => INIT_VAL_256,
      INIT_7B => INIT_VAL_256,
      INIT_7C => INIT_VAL_256,
      INIT_7D => INIT_VAL_256,
      INIT_7E => INIT_VAL_256,
      INIT_7F => INIT_VAL_256,
      INIT_A => INIT_VAL_36,
      INIT_B => INIT_VAL_36,
      INIT_FILE => string("NONE"),
      READ_WIDTH_A => 8,
      READ_WIDTH_B => 8,
      SIM_COLLISION_CHECK => "NONE",
      SIM_MODE => "SAFE",  -- This parameter is valid only for Virtex5
      SRVAL_A => INIT_VAL_36,
      SRVAL_B => INIT_VAL_36,
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B => "WRITE_FIRST",
      WRITE_WIDTH_A => 8,
      WRITE_WIDTH_B => 8,
      IS_CLKARDCLK_INVERTED  =>  '0',
      IS_CLKBWRCLK_INVERTED => '0',
      IS_ENARDEN_INVERTED => '0',
      IS_ENBWREN_INVERTED => '0',
      IS_RSTRAMARSTRAM_INVERTED => '0',
      IS_RSTRAMB_INVERTED => '0',
      IS_RSTREGARSTREG_INVERTED => '0',
      IS_RSTREGB_INVERTED => '0',
      RAM_EXTENSION_A =>  "NONE",
      RAM_EXTENSION_B => "NONE",
      RAM_MODE  => "TDP",
      RDADDR_COLLISION_HWCONFIG  =>  "DELAYED_WRITE",
      READ_WIDTH_A => 8,
      READ_WIDTH_B  => 0,
      RSTREG_PRIORITY_A  => "RSTREG",
      RSTREG_PRIORITY_B  => "RSTREG",
      SIM_COLLISION_CHECK  => "NONE", --"ALL",
      SIM_DEVICE  => "7SERIES",
      SRVAL_A  => INIT_VAL_36,
      SRVAL_B  => INIT_VAL_36,
      WRITE_MODE_A => "WRITE_FIRST",
      WRITE_MODE_B  => "WRITE_FIRST",
      WRITE_WIDTH_A  => 8,
      WRITE_WIDTH_B  => 8
    )
    port map (
      CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR  => open,
        DOADO => a_dout,
        DOBDO => b_dout,
        DOPADOP  => open,
        DOPBDOP  => open,
        ECCPARITY  => open,
        RDADDRECC  => open,
        SBITERR  => open,
        ADDRARDADDR => a_addr,
        ADDRBWRADDR => b_addr,
        CASCADEINA  => open,
        CASCADEINB  => open,
        CLKARDCLK => clka,
        CLKBWRCLK => clkb,
        DIADI => a_din,
      DIBDI => "00000000",
      DIPADIP => "0000",
      DIPBDIP => "0000",
      ENARDEN => '1',
      ENBWREN => '1',
      INJECTDBITERR => '0',
      INJECTSBITERR => '0',
      REGCEAREGCE => '0',
      REGCEB => '0',
      RSTRAMARSTRAM => '0',
      RSRSTRAMBTB => '0',
      RSTREGARSTREG => '0',
      RSTREGB => '0',
      WEA => data_we,
      WEBWE => '0'
      );
end arch;


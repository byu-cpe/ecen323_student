// Listing 13.1
// ROM with synchonous read (inferring Block RAM)
// character ROM
//   - 8-by-16 (8-by-2^4) font
//   - 128 (2^7) characters
//   - ROM size: 512-by-8 (2^11-by-8) bits
//               16K bits: 1 BRAM

module font_rom (
                 input logic clk,
                 input wire logic[10:0] addr,
                 output logic[7:0] data
                 );

   logic [10:0] addr_reg;
   logic [7:0]  rom[2048];

   initial begin
      rom[0] = 8'b00000000;  // 0
      rom[1] = 8'b00000000;  // 1
      rom[2] = 8'b00000000;  // 2
      rom[3] = 8'b00000000;  // 3
      rom[4] = 8'b00000000;  // 4
      rom[5] = 8'b00000000;  // 5
      rom[6] = 8'b00000000;  // 6
      rom[7] = 8'b00000000;  // 7
      rom[8] = 8'b00000000;  // 8
      rom[9] = 8'b00000000;  // 9
      rom[10] = 8'b00000000;  // a
      rom[11] = 8'b00000000;  // b
      rom[12] = 8'b00000000;  // c
      rom[13] = 8'b00000000;  // d
      rom[14] = 8'b00000000;  // e
      rom[15] = 8'b00000000;  // f
      // code x01
      rom[16] = 8'b00000000;  // 0
      rom[17] = 8'b00000000;  // 1
      rom[18] = 8'b01111110;  // 2  ******
      rom[19] = 8'b10000001;  // 3 *      *
      rom[20] = 8'b10100101;  // 4 * *  * *
      rom[21] = 8'b10000001;  // 5 *      *
      rom[22] = 8'b10000001;  // 6 *      *
      rom[23] = 8'b10111101;  // 7 * **** *
      rom[24] = 8'b10011001;  // 8 *  **  *
      rom[25] = 8'b10000001;  // 9 *      *
      rom[26] = 8'b10000001;  // a *      *
      rom[27] = 8'b01111110;  // b  ******
      rom[28] = 8'b00000000;  // c
      rom[29] = 8'b00000000;  // d
      rom[30] = 8'b00000000;  // e
      rom[31] = 8'b00000000;  // f
      // code x02
      rom[32] = 8'b00000000;  // 0
      rom[33] = 8'b00000000;  // 1
      rom[34] = 8'b01111110;  // 2  ******
      rom[35] = 8'b11111111;  // 3 ********
      rom[36] = 8'b11011011;  // 4 ** ** **
      rom[37] = 8'b11111111;  // 5 ********
      rom[38] = 8'b11111111;  // 6 ********
      rom[39] = 8'b11000011;  // 7 **    **
      rom[40] = 8'b11100111;  // 8 ***  ***
      rom[41] = 8'b11111111;  // 9 ********
      rom[42] = 8'b11111111;  // a ********
      rom[43] = 8'b01111110;  // b  ******
      rom[44] = 8'b00000000;  // c
      rom[45] = 8'b00000000;  // d
      rom[46] = 8'b00000000;  // e
      rom[47] = 8'b00000000;  // f
      // code x03
      rom[48] = 8'b00000000;  // 0
      rom[49] = 8'b00000000;  // 1
      rom[50] = 8'b00000000;  // 2
      rom[51] = 8'b00000000;  // 3
      rom[52] = 8'b01101100;  // 4  ** **
      rom[53] = 8'b11111110;  // 5 *******
      rom[54] = 8'b11111110;  // 6 *******
      rom[55] = 8'b11111110;  // 7 *******
      rom[56] = 8'b11111110;  // 8 *******
      rom[57] = 8'b01111100;  // 9  *****
      rom[58] = 8'b00111000;  // a   ***
      rom[59] = 8'b00010000;  // b    *
      rom[60] = 8'b00000000;  // c
      rom[61] = 8'b00000000;  // d
      rom[62] = 8'b00000000;  // e
      rom[63] = 8'b00000000;  // f
      // code x04
      rom[64] = 8'b00000000;  // 0
      rom[65] = 8'b00000000;  // 1
      rom[66] = 8'b00000000;  // 2
      rom[67] = 8'b00000000;  // 3
      rom[68] = 8'b00010000;  // 4    *
      rom[69] = 8'b00111000;  // 5   ***
      rom[70] = 8'b01111100;  // 6  *****
      rom[71] = 8'b11111110;  // 7 *******
      rom[72] = 8'b01111100;  // 8  *****
      rom[73] = 8'b00111000;  // 9   ***
      rom[74] = 8'b00010000;  // a    *
      rom[75] = 8'b00000000;  // b
      rom[76] = 8'b00000000;  // c
      rom[77] = 8'b00000000;  // d
      rom[78] = 8'b00000000;  // e
      rom[79] = 8'b00000000;  // f
      // code x05
      rom[80] = 8'b00000000;  // 0
      rom[81] = 8'b00000000;  // 1
      rom[82] = 8'b00000000;  // 2
      rom[83] = 8'b00011000;  // 3    **
      rom[84] = 8'b00111100;  // 4   ****
      rom[85] = 8'b00111100;  // 5   ****
      rom[86] = 8'b11100111;  // 6 ***  ***
      rom[87] = 8'b11100111;  // 7 ***  ***
      rom[88] = 8'b11100111;  // 8 ***  ***
      rom[89] = 8'b00011000;  // 9    **
      rom[90] = 8'b00011000;  // a    **
      rom[91] = 8'b00111100;  // b   ****
      rom[92] = 8'b00000000;  // c
      rom[93] = 8'b00000000;  // d
      rom[94] = 8'b00000000;  // e
      rom[95] = 8'b00000000;  // f
      // code x06
      rom[96] = 8'b00000000;  // 0
      rom[97] = 8'b00000000;  // 1
      rom[98] = 8'b00000000;  // 2
      rom[99] = 8'b00011000;  // 3    **
      rom[100] = 8'b00111100;  // 4   ****
      rom[101] = 8'b01111110;  // 5  ******
      rom[102] = 8'b11111111;  // 6 ********
      rom[103] = 8'b11111111;  // 7 ********
      rom[104] = 8'b01111110;  // 8  ******
      rom[105] = 8'b00011000;  // 9    **
      rom[106] = 8'b00011000;  // a    **
      rom[107] = 8'b00111100;  // b   ****
      rom[108] = 8'b00000000;  // c
      rom[109] = 8'b00000000;  // d
      rom[110] = 8'b00000000;  // e
      rom[111] = 8'b00000000;  // f
      // code x07
      rom[112] = 8'b00000000;  // 0
      rom[113] = 8'b00000000;  // 1
      rom[114] = 8'b00000000;  // 2
      rom[115] = 8'b00000000;  // 3
      rom[116] = 8'b00000000;  // 4
      rom[117] = 8'b00000000;  // 5
      rom[118] = 8'b00011000;  // 6    **
      rom[119] = 8'b00111100;  // 7   ****
      rom[120] = 8'b00111100;  // 8   ****
      rom[121] = 8'b00011000;  // 9    **
      rom[122] = 8'b00000000;  // a
      rom[123] = 8'b00000000;  // b
      rom[124] = 8'b00000000;  // c
      rom[125] = 8'b00000000;  // d
      rom[126] = 8'b00000000;  // e
      rom[127] = 8'b00000000;  // f
      // code x08
      rom[128] = 8'b11111111;  // 0 ********
      rom[129] = 8'b11111111;  // 1 ********
      rom[130] = 8'b11111111;  // 2 ********
      rom[131] = 8'b11111111;  // 3 ********
      rom[132] = 8'b11111111;  // 4 ********
      rom[133] = 8'b11111111;  // 5 ********
      rom[134] = 8'b11100111;  // 6 ***  ***
      rom[135] = 8'b11000011;  // 7 **    **
      rom[136] = 8'b11000011;  // 8 **    **
      rom[137] = 8'b11100111;  // 9 ***  ***
      rom[138] = 8'b11111111;  // a ********
      rom[139] = 8'b11111111;  // b ********
      rom[140] = 8'b11111111;  // c ********
      rom[141] = 8'b11111111;  // d ********
      rom[142] = 8'b11111111;  // e ********
      rom[143] = 8'b11111111;  // f ********
      // code x09
      rom[144] = 8'b00000000;  // 0
      rom[145] = 8'b00000000;  // 1
      rom[146] = 8'b00000000;  // 2
      rom[147] = 8'b00000000;  // 3
      rom[148] = 8'b00000000;  // 4
      rom[149] = 8'b00111100;  // 5   ****
      rom[150] = 8'b01100110;  // 6  **  **
      rom[151] = 8'b01000010;  // 7  *    *
      rom[152] = 8'b01000010;  // 8  *    *
      rom[153] = 8'b01100110;  // 9  **  **
      rom[154] = 8'b00111100;  // a   ****
      rom[155] = 8'b00000000;  // b
      rom[156] = 8'b00000000;  // c
      rom[157] = 8'b00000000;  // d
      rom[158] = 8'b00000000;  // e
      rom[159] = 8'b00000000;  // f
      // code x0a
      rom[160] = 8'b11111111;  // 0 ********
      rom[161] = 8'b11111111;  // 1 ********
      rom[162] = 8'b11111111;  // 2 ********
      rom[163] = 8'b11111111;  // 3 ********
      rom[164] = 8'b11111111;  // 4 ********
      rom[165] = 8'b11000011;  // 5 **    **
      rom[166] = 8'b10011001;  // 6 *  **  *
      rom[167] = 8'b10111101;  // 7 * **** *
      rom[168] = 8'b10111101;  // 8 * **** *
      rom[169] = 8'b10011001;  // 9 *  **  *
      rom[170] = 8'b11000011;  // a **    **
      rom[171] = 8'b11111111;  // b ********
      rom[172] = 8'b11111111;  // c ********
      rom[173] = 8'b11111111;  // d ********
      rom[174] = 8'b11111111;  // e ********
      rom[175] = 8'b11111111;  // f ********
      // code x0b
      rom[176] = 8'b00000000;  // 0
      rom[177] = 8'b00000000;  // 1
      rom[178] = 8'b00011110;  // 2    ****
      rom[179] = 8'b00001110;  // 3     ***
      rom[180] = 8'b00011010;  // 4    ** *
      rom[181] = 8'b00110010;  // 5   **  *
      rom[182] = 8'b01111000;  // 6  ****
      rom[183] = 8'b11001100;  // 7 **  **
      rom[184] = 8'b11001100;  // 8 **  **
      rom[185] = 8'b11001100;  // 9 **  **
      rom[186] = 8'b11001100;  // a **  **
      rom[187] = 8'b01111000;  // b  ****
      rom[188] = 8'b00000000;  // c
      rom[189] = 8'b00000000;  // d
      rom[190] = 8'b00000000;  // e
      rom[191] = 8'b00000000;  // f
      // code x0c
      rom[192] = 8'b00000000;  // 0
      rom[193] = 8'b00000000;  // 1
      rom[194] = 8'b00111100;  // 2   ****
      rom[195] = 8'b01100110;  // 3  **  **
      rom[196] = 8'b01100110;  // 4  **  **
      rom[197] = 8'b01100110;  // 5  **  **
      rom[198] = 8'b01100110;  // 6  **  **
      rom[199] = 8'b00111100;  // 7   ****
      rom[200] = 8'b00011000;  // 8    **
      rom[201] = 8'b01111110;  // 9  ******
      rom[202] = 8'b00011000;  // a    **
      rom[203] = 8'b00011000;  // b    **
      rom[204] = 8'b00000000;  // c
      rom[205] = 8'b00000000;  // d
      rom[206] = 8'b00000000;  // e
      rom[207] = 8'b00000000;  // f
      // code x0d
      rom[208] = 8'b00000000;  // 0
      rom[209] = 8'b00000000;  // 1
      rom[210] = 8'b00111111;  // 2   ******
      rom[211] = 8'b00110011;  // 3   **  **
      rom[212] = 8'b00111111;  // 4   ******
      rom[213] = 8'b00110000;  // 5   **
      rom[214] = 8'b00110000;  // 6   **
      rom[215] = 8'b00110000;  // 7   **
      rom[216] = 8'b00110000;  // 8   **
      rom[217] = 8'b01110000;  // 9  ***
      rom[218] = 8'b11110000;  // a ****
      rom[219] = 8'b11100000;  // b ***
      rom[220] = 8'b00000000;  // c
      rom[221] = 8'b00000000;  // d
      rom[222] = 8'b00000000;  // e
      rom[223] = 8'b00000000;  // f
      // code x0e
      rom[224] = 8'b00000000;  // 0
      rom[225] = 8'b00000000;  // 1
      rom[226] = 8'b01111111;  // 2  *******
      rom[227] = 8'b01100011;  // 3  **   **
      rom[228] = 8'b01111111;  // 4  *******
      rom[229] = 8'b01100011;  // 5  **   **
      rom[230] = 8'b01100011;  // 6  **   **
      rom[231] = 8'b01100011;  // 7  **   **
      rom[232] = 8'b01100011;  // 8  **   **
      rom[233] = 8'b01100111;  // 9  **  ***
      rom[234] = 8'b11100111;  // a ***  ***
      rom[235] = 8'b11100110;  // b ***  **
      rom[236] = 8'b11000000;  // c **
      rom[237] = 8'b00000000;  // d
      rom[238] = 8'b00000000;  // e
      rom[239] = 8'b00000000;  // f
      // code x0f
      rom[240] = 8'b00000000;  // 0
      rom[241] = 8'b00000000;  // 1
      rom[242] = 8'b00000000;  // 2
      rom[243] = 8'b00011000;  // 3    **
      rom[244] = 8'b00011000;  // 4    **
      rom[245] = 8'b11011011;  // 5 ** ** **
      rom[246] = 8'b00111100;  // 6   ****
      rom[247] = 8'b11100111;  // 7 ***  ***
      rom[248] = 8'b00111100;  // 8   ****
      rom[249] = 8'b11011011;  // 9 ** ** **
      rom[250] = 8'b00011000;  // a    **
      rom[251] = 8'b00011000;  // b    **
      rom[252] = 8'b00000000;  // c
      rom[253] = 8'b00000000;  // d
      rom[254] = 8'b00000000;  // e
      rom[255] = 8'b00000000;  // f
      // code x10
      rom[256] = 8'b00000000;  // 0
      rom[257] = 8'b10000000;  // 1 *
      rom[258] = 8'b11000000;  // 2 **
      rom[259] = 8'b11100000;  // 3 ***
      rom[260] = 8'b11110000;  // 4 ****
      rom[261] = 8'b11111000;  // 5 *****
      rom[262] = 8'b11111110;  // 6 *******
      rom[263] = 8'b11111000;  // 7 *****
      rom[264] = 8'b11110000;  // 8 ****
      rom[265] = 8'b11100000;  // 9 ***
      rom[266] = 8'b11000000;  // a **
      rom[267] = 8'b10000000;  // b *
      rom[268] = 8'b00000000;  // c
      rom[269] = 8'b00000000;  // d
      rom[270] = 8'b00000000;  // e
      rom[271] = 8'b00000000;  // f
      // code x11
      rom[272] = 8'b00000000;  // 0
      rom[273] = 8'b00000010;  // 1       *
      rom[274] = 8'b00000110;  // 2      **
      rom[275] = 8'b00001110;  // 3     ***
      rom[276] = 8'b00011110;  // 4    ****
      rom[277] = 8'b00111110;  // 5   *****
      rom[278] = 8'b11111110;  // 6 *******
      rom[279] = 8'b00111110;  // 7   *****
      rom[280] = 8'b00011110;  // 8    ****
      rom[281] = 8'b00001110;  // 9     ***
      rom[282] = 8'b00000110;  // a      **
      rom[283] = 8'b00000010;  // b       *
      rom[284] = 8'b00000000;  // c
      rom[285] = 8'b00000000;  // d
      rom[286] = 8'b00000000;  // e
      rom[287] = 8'b00000000;  // f
      // code x12
      rom[288] = 8'b00000000;  // 0
      rom[289] = 8'b00000000;  // 1
      rom[290] = 8'b00011000;  // 2    **
      rom[291] = 8'b00111100;  // 3   ****
      rom[292] = 8'b01111110;  // 4  ******
      rom[293] = 8'b00011000;  // 5    **
      rom[294] = 8'b00011000;  // 6    **
      rom[295] = 8'b00011000;  // 7    **
      rom[296] = 8'b01111110;  // 8  ******
      rom[297] = 8'b00111100;  // 9   ****
      rom[298] = 8'b00011000;  // a    **
      rom[299] = 8'b00000000;  // b
      rom[300] = 8'b00000000;  // c
      rom[301] = 8'b00000000;  // d
      rom[302] = 8'b00000000;  // e
      rom[303] = 8'b00000000;  // f
      // code x13
      rom[304] = 8'b00000000;  // 0
      rom[305] = 8'b00000000;  // 1
      rom[306] = 8'b01100110;  // 2  **  **
      rom[307] = 8'b01100110;  // 3  **  **
      rom[308] = 8'b01100110;  // 4  **  **
      rom[309] = 8'b01100110;  // 5  **  **
      rom[310] = 8'b01100110;  // 6  **  **
      rom[311] = 8'b01100110;  // 7  **  **
      rom[312] = 8'b01100110;  // 8  **  **
      rom[313] = 8'b00000000;  // 9
      rom[314] = 8'b01100110;  // a  **  **
      rom[315] = 8'b01100110;  // b  **  **
      rom[316] = 8'b00000000;  // c
      rom[317] = 8'b00000000;  // d
      rom[318] = 8'b00000000;  // e
      rom[319] = 8'b00000000;  // f
      // code x14
      rom[320] = 8'b00000000;  // 0
      rom[321] = 8'b00000000;  // 1
      rom[322] = 8'b01111111;  // 2  *******
      rom[323] = 8'b11011011;  // 3 ** ** **
      rom[324] = 8'b11011011;  // 4 ** ** **
      rom[325] = 8'b11011011;  // 5 ** ** **
      rom[326] = 8'b01111011;  // 6  **** **
      rom[327] = 8'b00011011;  // 7    ** **
      rom[328] = 8'b00011011;  // 8    ** **
      rom[329] = 8'b00011011;  // 9    ** **
      rom[330] = 8'b00011011;  // a    ** **
      rom[331] = 8'b00011011;  // b    ** **
      rom[332] = 8'b00000000;  // c
      rom[333] = 8'b00000000;  // d
      rom[334] = 8'b00000000;  // e
      rom[335] = 8'b00000000;  // f
      // code x15
      rom[336] = 8'b00000000;  // 0
      rom[337] = 8'b01111100;  // 1  *****
      rom[338] = 8'b11000110;  // 2 **   **
      rom[339] = 8'b01100000;  // 3  **
      rom[340] = 8'b00111000;  // 4   ***
      rom[341] = 8'b01101100;  // 5  ** **
      rom[342] = 8'b11000110;  // 6 **   **
      rom[343] = 8'b11000110;  // 7 **   **
      rom[344] = 8'b01101100;  // 8  ** **
      rom[345] = 8'b00111000;  // 9   ***
      rom[346] = 8'b00001100;  // a     **
      rom[347] = 8'b11000110;  // b **   **
      rom[348] = 8'b01111100;  // c  *****
      rom[349] = 8'b00000000;  // d
      rom[350] = 8'b00000000;  // e
      rom[351] = 8'b00000000;  // f
      // code x16
      rom[352] = 8'b00000000;  // 0
      rom[353] = 8'b00000000;  // 1
      rom[354] = 8'b00000000;  // 2
      rom[355] = 8'b00000000;  // 3
      rom[356] = 8'b00000000;  // 4
      rom[357] = 8'b00000000;  // 5
      rom[358] = 8'b00000000;  // 6
      rom[359] = 8'b00000000;  // 7
      rom[360] = 8'b11111110;  // 8 *******
      rom[361] = 8'b11111110;  // 9 *******
      rom[362] = 8'b11111110;  // a *******
      rom[363] = 8'b11111110;  // b *******
      rom[364] = 8'b00000000;  // c
      rom[365] = 8'b00000000;  // d
      rom[366] = 8'b00000000;  // e
      rom[367] = 8'b00000000;  // f
      // code x17
      rom[368] = 8'b00000000;  // 0
      rom[369] = 8'b00000000;  // 1
      rom[370] = 8'b00011000;  // 2    **
      rom[371] = 8'b00111100;  // 3   ****
      rom[372] = 8'b01111110;  // 4  ******
      rom[373] = 8'b00011000;  // 5    **
      rom[374] = 8'b00011000;  // 6    **
      rom[375] = 8'b00011000;  // 7    **
      rom[376] = 8'b01111110;  // 8  ******
      rom[377] = 8'b00111100;  // 9   ****
      rom[378] = 8'b00011000;  // a    **
      rom[379] = 8'b01111110;  // b  ******
      rom[380] = 8'b00110000;  // c
      rom[381] = 8'b00000000;  // d
      rom[382] = 8'b00000000;  // e
      rom[383] = 8'b00000000;  // f
      // code x18
      rom[384] = 8'b00000000;  // 0
      rom[385] = 8'b00000000;  // 1
      rom[386] = 8'b00011000;  // 2    **
      rom[387] = 8'b00111100;  // 3   ****
      rom[388] = 8'b01111110;  // 4  ******
      rom[389] = 8'b00011000;  // 5    **
      rom[390] = 8'b00011000;  // 6    **
      rom[391] = 8'b00011000;  // 7    **
      rom[392] = 8'b00011000;  // 8    **
      rom[393] = 8'b00011000;  // 9    **
      rom[394] = 8'b00011000;  // a    **
      rom[395] = 8'b00011000;  // b    **
      rom[396] = 8'b00000000;  // c
      rom[397] = 8'b00000000;  // d
      rom[398] = 8'b00000000;  // e
      rom[399] = 8'b00000000;  // f
      // code x19
      rom[400] = 8'b00000000;  // 0
      rom[401] = 8'b00000000;  // 1
      rom[402] = 8'b00011000;  // 2    **
      rom[403] = 8'b00011000;  // 3    **
      rom[404] = 8'b00011000;  // 4    **
      rom[405] = 8'b00011000;  // 5    **
      rom[406] = 8'b00011000;  // 6    **
      rom[407] = 8'b00011000;  // 7    **
      rom[408] = 8'b00011000;  // 8    **
      rom[409] = 8'b01111110;  // 9  ******
      rom[410] = 8'b00111100;  // a   ****
      rom[411] = 8'b00011000;  // b    **
      rom[412] = 8'b00000000;  // c
      rom[413] = 8'b00000000;  // d
      rom[414] = 8'b00000000;  // e
      rom[415] = 8'b00000000;  // f
      // code x1a
      rom[416] = 8'b00000000;  // 0
      rom[417] = 8'b00000000;  // 1
      rom[418] = 8'b00000000;  // 2
      rom[419] = 8'b00000000;  // 3
      rom[420] = 8'b00000000;  // 4
      rom[421] = 8'b00011000;  // 5    **
      rom[422] = 8'b00001100;  // 6     **
      rom[423] = 8'b11111110;  // 7 *******
      rom[424] = 8'b00001100;  // 8     **
      rom[425] = 8'b00011000;  // 9    **
      rom[426] = 8'b00000000;  // a
      rom[427] = 8'b00000000;  // b
      rom[428] = 8'b00000000;  // c
      rom[429] = 8'b00000000;  // d
      rom[430] = 8'b00000000;  // e
      rom[431] = 8'b00000000;  // f
      // code x1b
      rom[432] = 8'b00000000;  // 0
      rom[433] = 8'b00000000;  // 1
      rom[434] = 8'b00000000;  // 2
      rom[435] = 8'b00000000;  // 3
      rom[436] = 8'b00000000;  // 4
      rom[437] = 8'b00110000;  // 5   **
      rom[438] = 8'b01100000;  // 6  **
      rom[439] = 8'b11111110;  // 7 *******
      rom[440] = 8'b01100000;  // 8  **
      rom[441] = 8'b00110000;  // 9   **
      rom[442] = 8'b00000000;  // a
      rom[443] = 8'b00000000;  // b
      rom[444] = 8'b00000000;  // c
      rom[445] = 8'b00000000;  // d
      rom[446] = 8'b00000000;  // e
      rom[447] = 8'b00000000;  // f
      // code x1c
      rom[448] = 8'b00000000;  // 0
      rom[449] = 8'b00000000;  // 1
      rom[450] = 8'b00000000;  // 2
      rom[451] = 8'b00000000;  // 3
      rom[452] = 8'b00000000;  // 4
      rom[453] = 8'b00000000;  // 5
      rom[454] = 8'b11000000;  // 6 **
      rom[455] = 8'b11000000;  // 7 **
      rom[456] = 8'b11000000;  // 8 **
      rom[457] = 8'b11111110;  // 9 *******
      rom[458] = 8'b00000000;  // a
      rom[459] = 8'b00000000;  // b
      rom[460] = 8'b00000000;  // c
      rom[461] = 8'b00000000;  // d
      rom[462] = 8'b00000000;  // e
      rom[463] = 8'b00000000;  // f
      // code x1d
      rom[464] = 8'b00000000;  // 0
      rom[465] = 8'b00000000;  // 1
      rom[466] = 8'b00000000;  // 2
      rom[467] = 8'b00000000;  // 3
      rom[468] = 8'b00000000;  // 4
      rom[469] = 8'b00100100;  // 5   *  *
      rom[470] = 8'b01100110;  // 6  **  **
      rom[471] = 8'b11111111;  // 7 ********
      rom[472] = 8'b01100110;  // 8  **  **
      rom[473] = 8'b00100100;  // 9   *  *
      rom[474] = 8'b00000000;  // a
      rom[475] = 8'b00000000;  // b
      rom[476] = 8'b00000000;  // c
      rom[477] = 8'b00000000;  // d
      rom[478] = 8'b00000000;  // e
      rom[479] = 8'b00000000;  // f
      // code x1e
      rom[480] = 8'b00000000;  // 0
      rom[481] = 8'b00000000;  // 1
      rom[482] = 8'b00000000;  // 2
      rom[483] = 8'b00000000;  // 3
      rom[484] = 8'b00010000;  // 4    *
      rom[485] = 8'b00111000;  // 5   ***
      rom[486] = 8'b00111000;  // 6   ***
      rom[487] = 8'b01111100;  // 7  *****
      rom[488] = 8'b01111100;  // 8  *****
      rom[489] = 8'b11111110;  // 9 *******
      rom[490] = 8'b11111110;  // a *******
      rom[491] = 8'b00000000;  // b
      rom[492] = 8'b00000000;  // c
      rom[493] = 8'b00000000;  // d
      rom[494] = 8'b00000000;  // e
      rom[495] = 8'b00000000;  // f
      // code x1f
      rom[496] = 8'b00000000;  // 0
      rom[497] = 8'b00000000;  // 1
      rom[498] = 8'b00000000;  // 2
      rom[499] = 8'b00000000;  // 3
      rom[500] = 8'b11111110;  // 4 *******
      rom[501] = 8'b11111110;  // 5 *******
      rom[502] = 8'b01111100;  // 6  *****
      rom[503] = 8'b01111100;  // 7  *****
      rom[504] = 8'b00111000;  // 8   ***
      rom[505] = 8'b00111000;  // 9   ***
      rom[506] = 8'b00010000;  // a    *
      rom[507] = 8'b00000000;  // b
      rom[508] = 8'b00000000;  // c
      rom[509] = 8'b00000000;  // d
      rom[510] = 8'b00000000;  // e
      rom[511] = 8'b00000000;  // f
      // code x20
      rom[512] = 8'b00000000;  // 0
      rom[513] = 8'b00000000;  // 1
      rom[514] = 8'b00000000;  // 2
      rom[515] = 8'b00000000;  // 3
      rom[516] = 8'b00000000;  // 4
      rom[517] = 8'b00000000;  // 5
      rom[518] = 8'b00000000;  // 6
      rom[519] = 8'b00000000;  // 7
      rom[520] = 8'b00000000;  // 8
      rom[521] = 8'b00000000;  // 9
      rom[522] = 8'b00000000;  // a
      rom[523] = 8'b00000000;  // b
      rom[524] = 8'b00000000;  // c
      rom[525] = 8'b00000000;  // d
      rom[526] = 8'b00000000;  // e
      rom[527] = 8'b00000000;  // f
      // code x21
      rom[528] = 8'b00000000;  // 0
      rom[529] = 8'b00000000;  // 1
      rom[530] = 8'b00011000;  // 2    **
      rom[531] = 8'b00111100;  // 3   ****
      rom[532] = 8'b00111100;  // 4   ****
      rom[533] = 8'b00111100;  // 5   ****
      rom[534] = 8'b00011000;  // 6    **
      rom[535] = 8'b00011000;  // 7    **
      rom[536] = 8'b00011000;  // 8    **
      rom[537] = 8'b00000000;  // 9
      rom[538] = 8'b00011000;  // a    **
      rom[539] = 8'b00011000;  // b    **
      rom[540] = 8'b00000000;  // c
      rom[541] = 8'b00000000;  // d
      rom[542] = 8'b00000000;  // e
      rom[543] = 8'b00000000;  // f
      // code x22
      rom[544] = 8'b00000000;  // 0
      rom[545] = 8'b01100110;  // 1  **  **
      rom[546] = 8'b01100110;  // 2  **  **
      rom[547] = 8'b01100110;  // 3  **  **
      rom[548] = 8'b00100100;  // 4   *  *
      rom[549] = 8'b00000000;  // 5
      rom[550] = 8'b00000000;  // 6
      rom[551] = 8'b00000000;  // 7
      rom[552] = 8'b00000000;  // 8
      rom[553] = 8'b00000000;  // 9
      rom[554] = 8'b00000000;  // a
      rom[555] = 8'b00000000;  // b
      rom[556] = 8'b00000000;  // c
      rom[557] = 8'b00000000;  // d
      rom[558] = 8'b00000000;  // e
      rom[559] = 8'b00000000;  // f
      // code x23
      rom[560] = 8'b00000000;  // 0
      rom[561] = 8'b00000000;  // 1
      rom[562] = 8'b00000000;  // 2
      rom[563] = 8'b01101100;  // 3  ** **
      rom[564] = 8'b01101100;  // 4  ** **
      rom[565] = 8'b11111110;  // 5 *******
      rom[566] = 8'b01101100;  // 6  ** **
      rom[567] = 8'b01101100;  // 7  ** **
      rom[568] = 8'b01101100;  // 8  ** **
      rom[569] = 8'b11111110;  // 9 *******
      rom[570] = 8'b01101100;  // a  ** **
      rom[571] = 8'b01101100;  // b  ** **
      rom[572] = 8'b00000000;  // c
      rom[573] = 8'b00000000;  // d
      rom[574] = 8'b00000000;  // e
      rom[575] = 8'b00000000;  // f
      // code x24
      rom[576] = 8'b00011000;  // 0     **
      rom[577] = 8'b00011000;  // 1     **
      rom[578] = 8'b01111100;  // 2   *****
      rom[579] = 8'b11000110;  // 3  **   **
      rom[580] = 8'b11000010;  // 4  **    *
      rom[581] = 8'b11000000;  // 5  **
      rom[582] = 8'b01111100;  // 6   *****
      rom[583] = 8'b00000110;  // 7       **
      rom[584] = 8'b00000110;  // 8       **
      rom[585] = 8'b10000110;  // 9  *    **
      rom[586] = 8'b11000110;  // a  **   **
      rom[587] = 8'b01111100;  // b   *****
      rom[588] = 8'b00011000;  // c     **
      rom[589] = 8'b00011000;  // d     **
      rom[590] = 8'b00000000;  // e
      rom[591] = 8'b00000000;  // f
      // code x25
      rom[592] = 8'b00000000;  // 0
      rom[593] = 8'b00000000;  // 1
      rom[594] = 8'b00000000;  // 2
      rom[595] = 8'b00000000;  // 3
      rom[596] = 8'b11000010;  // 4 **    *
      rom[597] = 8'b11000110;  // 5 **   **
      rom[598] = 8'b00001100;  // 6     **
      rom[599] = 8'b00011000;  // 7    **
      rom[600] = 8'b00110000;  // 8   **
      rom[601] = 8'b01100000;  // 9  **
      rom[602] = 8'b11000110;  // a **   **
      rom[603] = 8'b10000110;  // b *    **
      rom[604] = 8'b00000000;  // c
      rom[605] = 8'b00000000;  // d
      rom[606] = 8'b00000000;  // e
      rom[607] = 8'b00000000;  // f
      // code x26
      rom[608] = 8'b00000000;  // 0
      rom[609] = 8'b00000000;  // 1
      rom[610] = 8'b00111000;  // 2   ***
      rom[611] = 8'b01101100;  // 3  ** **
      rom[612] = 8'b01101100;  // 4  ** **
      rom[613] = 8'b00111000;  // 5   ***
      rom[614] = 8'b01110110;  // 6  *** **
      rom[615] = 8'b11011100;  // 7 ** ***
      rom[616] = 8'b11001100;  // 8 **  **
      rom[617] = 8'b11001100;  // 9 **  **
      rom[618] = 8'b11001100;  // a **  **
      rom[619] = 8'b01110110;  // b  *** **
      rom[620] = 8'b00000000;  // c
      rom[621] = 8'b00000000;  // d
      rom[622] = 8'b00000000;  // e
      rom[623] = 8'b00000000;  // f
      // code x27
      rom[624] = 8'b00000000;  // 0
      rom[625] = 8'b00110000;  // 1   **
      rom[626] = 8'b00110000;  // 2   **
      rom[627] = 8'b00110000;  // 3   **
      rom[628] = 8'b01100000;  // 4  **
      rom[629] = 8'b00000000;  // 5
      rom[630] = 8'b00000000;  // 6
      rom[631] = 8'b00000000;  // 7
      rom[632] = 8'b00000000;  // 8
      rom[633] = 8'b00000000;  // 9
      rom[634] = 8'b00000000;  // a
      rom[635] = 8'b00000000;  // b
      rom[636] = 8'b00000000;  // c
      rom[637] = 8'b00000000;  // d
      rom[638] = 8'b00000000;  // e
      rom[639] = 8'b00000000;  // f
      // code x28
      rom[640] = 8'b00000000;  // 0
      rom[641] = 8'b00000000;  // 1
      rom[642] = 8'b00001100;  // 2     **
      rom[643] = 8'b00011000;  // 3    **
      rom[644] = 8'b00110000;  // 4   **
      rom[645] = 8'b00110000;  // 5   **
      rom[646] = 8'b00110000;  // 6   **
      rom[647] = 8'b00110000;  // 7   **
      rom[648] = 8'b00110000;  // 8   **
      rom[649] = 8'b00110000;  // 9   **
      rom[650] = 8'b00011000;  // a    **
      rom[651] = 8'b00001100;  // b     **
      rom[652] = 8'b00000000;  // c
      rom[653] = 8'b00000000;  // d
      rom[654] = 8'b00000000;  // e
      rom[655] = 8'b00000000;  // f
      // code x29
      rom[656] = 8'b00000000;  // 0
      rom[657] = 8'b00000000;  // 1
      rom[658] = 8'b00110000;  // 2   **
      rom[659] = 8'b00011000;  // 3    **
      rom[660] = 8'b00001100;  // 4     **
      rom[661] = 8'b00001100;  // 5     **
      rom[662] = 8'b00001100;  // 6     **
      rom[663] = 8'b00001100;  // 7     **
      rom[664] = 8'b00001100;  // 8     **
      rom[665] = 8'b00001100;  // 9     **
      rom[666] = 8'b00011000;  // a    **
      rom[667] = 8'b00110000;  // b   **
      rom[668] = 8'b00000000;  // c
      rom[669] = 8'b00000000;  // d
      rom[670] = 8'b00000000;  // e
      rom[671] = 8'b00000000;  // f
      // code x2a
      rom[672] = 8'b00000000;  // 0
      rom[673] = 8'b00000000;  // 1
      rom[674] = 8'b00000000;  // 2
      rom[675] = 8'b00000000;  // 3
      rom[676] = 8'b00000000;  // 4
      rom[677] = 8'b01100110;  // 5  **  **
      rom[678] = 8'b00111100;  // 6   ****
      rom[679] = 8'b11111111;  // 7 ********
      rom[680] = 8'b00111100;  // 8   ****
      rom[681] = 8'b01100110;  // 9  **  **
      rom[682] = 8'b00000000;  // a
      rom[683] = 8'b00000000;  // b
      rom[684] = 8'b00000000;  // c
      rom[685] = 8'b00000000;  // d
      rom[686] = 8'b00000000;  // e
      rom[687] = 8'b00000000;  // f
      // code x2b
      rom[688] = 8'b00000000;  // 0
      rom[689] = 8'b00000000;  // 1
      rom[690] = 8'b00000000;  // 2
      rom[691] = 8'b00000000;  // 3
      rom[692] = 8'b00000000;  // 4
      rom[693] = 8'b00011000;  // 5    **
      rom[694] = 8'b00011000;  // 6    **
      rom[695] = 8'b01111110;  // 7  ******
      rom[696] = 8'b00011000;  // 8    **
      rom[697] = 8'b00011000;  // 9    **
      rom[698] = 8'b00000000;  // a
      rom[699] = 8'b00000000;  // b
      rom[700] = 8'b00000000;  // c
      rom[701] = 8'b00000000;  // d
      rom[702] = 8'b00000000;  // e
      rom[703] = 8'b00000000;  // f
      // code x2c
      rom[704] = 8'b00000000;  // 0
      rom[705] = 8'b00000000;  // 1
      rom[706] = 8'b00000000;  // 2
      rom[707] = 8'b00000000;  // 3
      rom[708] = 8'b00000000;  // 4
      rom[709] = 8'b00000000;  // 5
      rom[710] = 8'b00000000;  // 6
      rom[711] = 8'b00000000;  // 7
      rom[712] = 8'b00000000;  // 8
      rom[713] = 8'b00011000;  // 9    **
      rom[714] = 8'b00011000;  // a    **
      rom[715] = 8'b00011000;  // b    **
      rom[716] = 8'b00110000;  // c   **
      rom[717] = 8'b00000000;  // d
      rom[718] = 8'b00000000;  // e
      rom[719] = 8'b00000000;  // f
      // code x2d
      rom[720] = 8'b00000000;  // 0
      rom[721] = 8'b00000000;  // 1
      rom[722] = 8'b00000000;  // 2
      rom[723] = 8'b00000000;  // 3
      rom[724] = 8'b00000000;  // 4
      rom[725] = 8'b00000000;  // 5
      rom[726] = 8'b00000000;  // 6
      rom[727] = 8'b01111110;  // 7  ******
      rom[728] = 8'b00000000;  // 8
      rom[729] = 8'b00000000;  // 9
      rom[730] = 8'b00000000;  // a
      rom[731] = 8'b00000000;  // b
      rom[732] = 8'b00000000;  // c
      rom[733] = 8'b00000000;  // d
      rom[734] = 8'b00000000;  // e
      rom[735] = 8'b00000000;  // f
      // code x2e
      rom[736] = 8'b00000000;  // 0
      rom[737] = 8'b00000000;  // 1
      rom[738] = 8'b00000000;  // 2
      rom[739] = 8'b00000000;  // 3
      rom[740] = 8'b00000000;  // 4
      rom[741] = 8'b00000000;  // 5
      rom[742] = 8'b00000000;  // 6
      rom[743] = 8'b00000000;  // 7
      rom[744] = 8'b00000000;  // 8
      rom[745] = 8'b00000000;  // 9
      rom[746] = 8'b00011000;  // a    **
      rom[747] = 8'b00011000;  // b    **
      rom[748] = 8'b00000000;  // c
      rom[749] = 8'b00000000;  // d
      rom[750] = 8'b00000000;  // e
      rom[751] = 8'b00000000;  // f
      // code x2f
      rom[752] = 8'b00000000;  // 0
      rom[753] = 8'b00000000;  // 1
      rom[754] = 8'b00000000;  // 2
      rom[755] = 8'b00000000;  // 3
      rom[756] = 8'b00000010;  // 4       *
      rom[757] = 8'b00000110;  // 5      **
      rom[758] = 8'b00001100;  // 6     **
      rom[759] = 8'b00011000;  // 7    **
      rom[760] = 8'b00110000;  // 8   **
      rom[761] = 8'b01100000;  // 9  **
      rom[762] = 8'b11000000;  // a **
      rom[763] = 8'b10000000;  // b *
      rom[764] = 8'b00000000;  // c
      rom[765] = 8'b00000000;  // d
      rom[766] = 8'b00000000;  // e
      rom[767] = 8'b00000000;  // f
      // code x30
      rom[768] = 8'b00000000;  // 0
      rom[769] = 8'b00000000;  // 1
      rom[770] = 8'b01111100;  // 2  *****
      rom[771] = 8'b11000110;  // 3 **   **
      rom[772] = 8'b11000110;  // 4 **   **
      rom[773] = 8'b11001110;  // 5 **  ***
      rom[774] = 8'b11011110;  // 6 ** ****
      rom[775] = 8'b11110110;  // 7 **** **
      rom[776] = 8'b11100110;  // 8 ***  **
      rom[777] = 8'b11000110;  // 9 **   **
      rom[778] = 8'b11000110;  // a **   **
      rom[779] = 8'b01111100;  // b  *****
      rom[780] = 8'b00000000;  // c
      rom[781] = 8'b00000000;  // d
      rom[782] = 8'b00000000;  // e
      rom[783] = 8'b00000000;  // f
      // code x31
      rom[784] = 8'b00000000;  // 0
      rom[785] = 8'b00000000;  // 1
      rom[786] = 8'b00011000;  // 2
      rom[787] = 8'b00111000;  // 3
      rom[788] = 8'b01111000;  // 4    **
      rom[789] = 8'b00011000;  // 5   ***
      rom[790] = 8'b00011000;  // 6  ****
      rom[791] = 8'b00011000;  // 7    **
      rom[792] = 8'b00011000;  // 8    **
      rom[793] = 8'b00011000;  // 9    **
      rom[794] = 8'b00011000;  // a    **
      rom[795] = 8'b01111110;  // b    **
      rom[796] = 8'b00000000;  // c    **
      rom[797] = 8'b00000000;  // d  ******
      rom[798] = 8'b00000000;  // e
      rom[799] = 8'b00000000;  // f
      // code x32
      rom[800] = 8'b00000000;  // 0
      rom[801] = 8'b00000000;  // 1
      rom[802] = 8'b01111100;  // 2  *****
      rom[803] = 8'b11000110;  // 3 **   **
      rom[804] = 8'b00000110;  // 4      **
      rom[805] = 8'b00001100;  // 5     **
      rom[806] = 8'b00011000;  // 6    **
      rom[807] = 8'b00110000;  // 7   **
      rom[808] = 8'b01100000;  // 8  **
      rom[809] = 8'b11000000;  // 9 **
      rom[810] = 8'b11000110;  // a **   **
      rom[811] = 8'b11111110;  // b *******
      rom[812] = 8'b00000000;  // c
      rom[813] = 8'b00000000;  // d
      rom[814] = 8'b00000000;  // e
      rom[815] = 8'b00000000;  // f
      // code x33
      rom[816] = 8'b00000000;  // 0
      rom[817] = 8'b00000000;  // 1
      rom[818] = 8'b01111100;  // 2  *****
      rom[819] = 8'b11000110;  // 3 **   **
      rom[820] = 8'b00000110;  // 4      **
      rom[821] = 8'b00000110;  // 5      **
      rom[822] = 8'b00111100;  // 6   ****
      rom[823] = 8'b00000110;  // 7      **
      rom[824] = 8'b00000110;  // 8      **
      rom[825] = 8'b00000110;  // 9      **
      rom[826] = 8'b11000110;  // a **   **
      rom[827] = 8'b01111100;  // b  *****
      rom[828] = 8'b00000000;  // c
      rom[829] = 8'b00000000;  // d
      rom[830] = 8'b00000000;  // e
      rom[831] = 8'b00000000;  // f
      // code x34
      rom[832] = 8'b00000000;  // 0
      rom[833] = 8'b00000000;  // 1
      rom[834] = 8'b00001100;  // 2     **
      rom[835] = 8'b00011100;  // 3    ***
      rom[836] = 8'b00111100;  // 4   ****
      rom[837] = 8'b01101100;  // 5  ** **
      rom[838] = 8'b11001100;  // 6 **  **
      rom[839] = 8'b11111110;  // 7 *******
      rom[840] = 8'b00001100;  // 8     **
      rom[841] = 8'b00001100;  // 9     **
      rom[842] = 8'b00001100;  // a     **
      rom[843] = 8'b00011110;  // b    ****
      rom[844] = 8'b00000000;  // c
      rom[845] = 8'b00000000;  // d
      rom[846] = 8'b00000000;  // e
      rom[847] = 8'b00000000;  // f
      // code x35
      rom[848] = 8'b00000000;  // 0
      rom[849] = 8'b00000000;  // 1
      rom[850] = 8'b11111110;  // 2 *******
      rom[851] = 8'b11000000;  // 3 **
      rom[852] = 8'b11000000;  // 4 **
      rom[853] = 8'b11000000;  // 5 **
      rom[854] = 8'b11111100;  // 6 ******
      rom[855] = 8'b00000110;  // 7      **
      rom[856] = 8'b00000110;  // 8      **
      rom[857] = 8'b00000110;  // 9      **
      rom[858] = 8'b11000110;  // a **   **
      rom[859] = 8'b01111100;  // b  *****
      rom[860] = 8'b00000000;  // c
      rom[861] = 8'b00000000;  // d
      rom[862] = 8'b00000000;  // e
      rom[863] = 8'b00000000;  // f
      // code x36
      rom[864] = 8'b00000000;  // 0
      rom[865] = 8'b00000000;  // 1
      rom[866] = 8'b00111000;  // 2   ***
      rom[867] = 8'b01100000;  // 3  **
      rom[868] = 8'b11000000;  // 4 **
      rom[869] = 8'b11000000;  // 5 **
      rom[870] = 8'b11111100;  // 6 ******
      rom[871] = 8'b11000110;  // 7 **   **
      rom[872] = 8'b11000110;  // 8 **   **
      rom[873] = 8'b11000110;  // 9 **   **
      rom[874] = 8'b11000110;  // a **   **
      rom[875] = 8'b01111100;  // b  *****
      rom[876] = 8'b00000000;  // c
      rom[877] = 8'b00000000;  // d
      rom[878] = 8'b00000000;  // e
      rom[879] = 8'b00000000;  // f
      // code x37
      rom[880] = 8'b00000000;  // 0
      rom[881] = 8'b00000000;  // 1
      rom[882] = 8'b11111110;  // 2 *******
      rom[883] = 8'b11000110;  // 3 **   **
      rom[884] = 8'b00000110;  // 4      **
      rom[885] = 8'b00000110;  // 5      **
      rom[886] = 8'b00001100;  // 6     **
      rom[887] = 8'b00011000;  // 7    **
      rom[888] = 8'b00110000;  // 8   **
      rom[889] = 8'b00110000;  // 9   **
      rom[890] = 8'b00110000;  // a   **
      rom[891] = 8'b00110000;  // b   **
      rom[892] = 8'b00000000;  // c
      rom[893] = 8'b00000000;  // d
      rom[894] = 8'b00000000;  // e
      rom[895] = 8'b00000000;  // f
      // code x38
      rom[896] = 8'b00000000;  // 0
      rom[897] = 8'b00000000;  // 1
      rom[898] = 8'b01111100;  // 2  *****
      rom[899] = 8'b11000110;  // 3 **   **
      rom[900] = 8'b11000110;  // 4 **   **
      rom[901] = 8'b11000110;  // 5 **   **
      rom[902] = 8'b01111100;  // 6  *****
      rom[903] = 8'b11000110;  // 7 **   **
      rom[904] = 8'b11000110;  // 8 **   **
      rom[905] = 8'b11000110;  // 9 **   **
      rom[906] = 8'b11000110;  // a **   **
      rom[907] = 8'b01111100;  // b  *****
      rom[908] = 8'b00000000;  // c
      rom[909] = 8'b00000000;  // d
      rom[910] = 8'b00000000;  // e
      rom[911] = 8'b00000000;  // f
      // code x39
      rom[912] = 8'b00000000;  // 0
      rom[913] = 8'b00000000;  // 1
      rom[914] = 8'b01111100;  // 2  *****
      rom[915] = 8'b11000110;  // 3 **   **
      rom[916] = 8'b11000110;  // 4 **   **
      rom[917] = 8'b11000110;  // 5 **   **
      rom[918] = 8'b01111110;  // 6  ******
      rom[919] = 8'b00000110;  // 7      **
      rom[920] = 8'b00000110;  // 8      **
      rom[921] = 8'b00000110;  // 9      **
      rom[922] = 8'b00001100;  // a     **
      rom[923] = 8'b01111000;  // b  ****
      rom[924] = 8'b00000000;  // c
      rom[925] = 8'b00000000;  // d
      rom[926] = 8'b00000000;  // e
      rom[927] = 8'b00000000;  // f
      // code x3a
      rom[928] = 8'b00000000;  // 0
      rom[929] = 8'b00000000;  // 1
      rom[930] = 8'b00000000;  // 2
      rom[931] = 8'b00000000;  // 3
      rom[932] = 8'b00011000;  // 4    **
      rom[933] = 8'b00011000;  // 5    **
      rom[934] = 8'b00000000;  // 6
      rom[935] = 8'b00000000;  // 7
      rom[936] = 8'b00000000;  // 8
      rom[937] = 8'b00011000;  // 9    **
      rom[938] = 8'b00011000;  // a    **
      rom[939] = 8'b00000000;  // b
      rom[940] = 8'b00000000;  // c
      rom[941] = 8'b00000000;  // d
      rom[942] = 8'b00000000;  // e
      rom[943] = 8'b00000000;  // f
      // code x3b
      rom[944] = 8'b00000000;  // 0
      rom[945] = 8'b00000000;  // 1
      rom[946] = 8'b00000000;  // 2
      rom[947] = 8'b00000000;  // 3
      rom[948] = 8'b00011000;  // 4    **
      rom[949] = 8'b00011000;  // 5    **
      rom[950] = 8'b00000000;  // 6
      rom[951] = 8'b00000000;  // 7
      rom[952] = 8'b00000000;  // 8
      rom[953] = 8'b00011000;  // 9    **
      rom[954] = 8'b00011000;  // a    **
      rom[955] = 8'b00110000;  // b   **
      rom[956] = 8'b00000000;  // c
      rom[957] = 8'b00000000;  // d
      rom[958] = 8'b00000000;  // e
      rom[959] = 8'b00000000;  // f
      // code x3c
      rom[960] = 8'b00000000;  // 0
      rom[961] = 8'b00000000;  // 1
      rom[962] = 8'b00000000;  // 2
      rom[963] = 8'b00000110;  // 3      **
      rom[964] = 8'b00001100;  // 4     **
      rom[965] = 8'b00011000;  // 5    **
      rom[966] = 8'b00110000;  // 6   **
      rom[967] = 8'b01100000;  // 7  **
      rom[968] = 8'b00110000;  // 8   **
      rom[969] = 8'b00011000;  // 9    **
      rom[970] = 8'b00001100;  // a     **
      rom[971] = 8'b00000110;  // b      **
      rom[972] = 8'b00000000;  // c
      rom[973] = 8'b00000000;  // d
      rom[974] = 8'b00000000;  // e
      rom[975] = 8'b00000000;  // f
      // code x3d
      rom[976] = 8'b00000000;  // 0
      rom[977] = 8'b00000000;  // 1
      rom[978] = 8'b00000000;  // 2
      rom[979] = 8'b00000000;  // 3
      rom[980] = 8'b00000000;  // 4
      rom[981] = 8'b01111110;  // 5  ******
      rom[982] = 8'b00000000;  // 6
      rom[983] = 8'b00000000;  // 7
      rom[984] = 8'b01111110;  // 8  ******
      rom[985] = 8'b00000000;  // 9
      rom[986] = 8'b00000000;  // a
      rom[987] = 8'b00000000;  // b
      rom[988] = 8'b00000000;  // c
      rom[989] = 8'b00000000;  // d
      rom[990] = 8'b00000000;  // e
      rom[991] = 8'b00000000;  // f
      // code x3e
      rom[992] = 8'b00000000;  // 0
      rom[993] = 8'b00000000;  // 1
      rom[994] = 8'b00000000;  // 2
      rom[995] = 8'b01100000;  // 3  **
      rom[996] = 8'b00110000;  // 4   **
      rom[997] = 8'b00011000;  // 5    **
      rom[998] = 8'b00001100;  // 6     **
      rom[999] = 8'b00000110;  // 7      **
      rom[1000] = 8'b00001100;  // 8     **
      rom[1001] = 8'b00011000;  // 9    **
      rom[1002] = 8'b00110000;  // a   **
      rom[1003] = 8'b01100000;  // b  **
      rom[1004] = 8'b00000000;  // c
      rom[1005] = 8'b00000000;  // d
      rom[1006] = 8'b00000000;  // e
      rom[1007] = 8'b00000000;  // f
      // code x3f
      rom[1008] = 8'b00000000;  // 0
      rom[1009] = 8'b00000000;  // 1
      rom[1010] = 8'b01111100;  // 2  *****
      rom[1011] = 8'b11000110;  // 3 **   **
      rom[1012] = 8'b11000110;  // 4 **   **
      rom[1013] = 8'b00001100;  // 5     **
      rom[1014] = 8'b00011000;  // 6    **
      rom[1015] = 8'b00011000;  // 7    **
      rom[1016] = 8'b00011000;  // 8    **
      rom[1017] = 8'b00000000;  // 9
      rom[1018] = 8'b00011000;  // a    **
      rom[1019] = 8'b00011000;  // b    **
      rom[1020] = 8'b00000000;  // c
      rom[1021] = 8'b00000000;  // d
      rom[1022] = 8'b00000000;  // e
      rom[1023] = 8'b00000000;  // f
      // code x40
      rom[1024] = 8'b00000000;  // 0
      rom[1025] = 8'b00000000;  // 1
      rom[1026] = 8'b01111100;  // 2  *****
      rom[1027] = 8'b11000110;  // 3 **   **
      rom[1028] = 8'b11000110;  // 4 **   **
      rom[1029] = 8'b11000110;  // 5 **   **
      rom[1030] = 8'b11011110;  // 6 ** ****
      rom[1031] = 8'b11011110;  // 7 ** ****
      rom[1032] = 8'b11011110;  // 8 ** ****
      rom[1033] = 8'b11011100;  // 9 ** ***
      rom[1034] = 8'b11000000;  // a **
      rom[1035] = 8'b01111100;  // b  *****
      rom[1036] = 8'b00000000;  // c
      rom[1037] = 8'b00000000;  // d
      rom[1038] = 8'b00000000;  // e
      rom[1039] = 8'b00000000;  // f
      // code x41
      rom[1040] = 8'b00000000;  // 0
      rom[1041] = 8'b00000000;  // 1
      rom[1042] = 8'b00010000;  // 2    *
      rom[1043] = 8'b00111000;  // 3   ***
      rom[1044] = 8'b01101100;  // 4  ** **
      rom[1045] = 8'b11000110;  // 5 **   **
      rom[1046] = 8'b11000110;  // 6 **   **
      rom[1047] = 8'b11111110;  // 7 *******
      rom[1048] = 8'b11000110;  // 8 **   **
      rom[1049] = 8'b11000110;  // 9 **   **
      rom[1050] = 8'b11000110;  // a **   **
      rom[1051] = 8'b11000110;  // b **   **
      rom[1052] = 8'b00000000;  // c
      rom[1053] = 8'b00000000;  // d
      rom[1054] = 8'b00000000;  // e
      rom[1055] = 8'b00000000;  // f
      // code x42
      rom[1056] = 8'b00000000;  // 0
      rom[1057] = 8'b00000000;  // 1
      rom[1058] = 8'b11111100;  // 2 ******
      rom[1059] = 8'b01100110;  // 3  **  **
      rom[1060] = 8'b01100110;  // 4  **  **
      rom[1061] = 8'b01100110;  // 5  **  **
      rom[1062] = 8'b01111100;  // 6  *****
      rom[1063] = 8'b01100110;  // 7  **  **
      rom[1064] = 8'b01100110;  // 8  **  **
      rom[1065] = 8'b01100110;  // 9  **  **
      rom[1066] = 8'b01100110;  // a  **  **
      rom[1067] = 8'b11111100;  // b ******
      rom[1068] = 8'b00000000;  // c
      rom[1069] = 8'b00000000;  // d
      rom[1070] = 8'b00000000;  // e
      rom[1071] = 8'b00000000;  // f
      // code x43
      rom[1072] = 8'b00000000;  // 0
      rom[1073] = 8'b00000000;  // 1
      rom[1074] = 8'b00111100;  // 2   ****
      rom[1075] = 8'b01100110;  // 3  **  **
      rom[1076] = 8'b11000010;  // 4 **    *
      rom[1077] = 8'b11000000;  // 5 **
      rom[1078] = 8'b11000000;  // 6 **
      rom[1079] = 8'b11000000;  // 7 **
      rom[1080] = 8'b11000000;  // 8 **
      rom[1081] = 8'b11000010;  // 9 **    *
      rom[1082] = 8'b01100110;  // a  **  **
      rom[1083] = 8'b00111100;  // b   ****
      rom[1084] = 8'b00000000;  // c
      rom[1085] = 8'b00000000;  // d
      rom[1086] = 8'b00000000;  // e
      rom[1087] = 8'b00000000;  // f
      // code x44
      rom[1088] = 8'b00000000;  // 0
      rom[1089] = 8'b00000000;  // 1
      rom[1090] = 8'b11111000;  // 2 *****
      rom[1091] = 8'b01101100;  // 3  ** **
      rom[1092] = 8'b01100110;  // 4  **  **
      rom[1093] = 8'b01100110;  // 5  **  **
      rom[1094] = 8'b01100110;  // 6  **  **
      rom[1095] = 8'b01100110;  // 7  **  **
      rom[1096] = 8'b01100110;  // 8  **  **
      rom[1097] = 8'b01100110;  // 9  **  **
      rom[1098] = 8'b01101100;  // a  ** **
      rom[1099] = 8'b11111000;  // b *****
      rom[1100] = 8'b00000000;  // c
      rom[1101] = 8'b00000000;  // d
      rom[1102] = 8'b00000000;  // e
      rom[1103] = 8'b00000000;  // f
      // code x45
      rom[1104] = 8'b00000000;  // 0
      rom[1105] = 8'b00000000;  // 1
      rom[1106] = 8'b11111110;  // 2 *******
      rom[1107] = 8'b01100110;  // 3  **  **
      rom[1108] = 8'b01100010;  // 4  **   *
      rom[1109] = 8'b01101000;  // 5  ** *
      rom[1110] = 8'b01111000;  // 6  ****
      rom[1111] = 8'b01101000;  // 7  ** *
      rom[1112] = 8'b01100000;  // 8  **
      rom[1113] = 8'b01100010;  // 9  **   *
      rom[1114] = 8'b01100110;  // a  **  **
      rom[1115] = 8'b11111110;  // b *******
      rom[1116] = 8'b00000000;  // c
      rom[1117] = 8'b00000000;  // d
      rom[1118] = 8'b00000000;  // e
      rom[1119] = 8'b00000000;  // f
      // code x46
      rom[1120] = 8'b00000000;  // 0
      rom[1121] = 8'b00000000;  // 1
      rom[1122] = 8'b11111110;  // 2 *******
      rom[1123] = 8'b01100110;  // 3  **  **
      rom[1124] = 8'b01100010;  // 4  **   *
      rom[1125] = 8'b01101000;  // 5  ** *
      rom[1126] = 8'b01111000;  // 6  ****
      rom[1127] = 8'b01101000;  // 7  ** *
      rom[1128] = 8'b01100000;  // 8  **
      rom[1129] = 8'b01100000;  // 9  **
      rom[1130] = 8'b01100000;  // a  **
      rom[1131] = 8'b11110000;  // b ****
      rom[1132] = 8'b00000000;  // c
      rom[1133] = 8'b00000000;  // d
      rom[1134] = 8'b00000000;  // e
      rom[1135] = 8'b00000000;  // f
      // code x47
      rom[1136] = 8'b00000000;  // 0
      rom[1137] = 8'b00000000;  // 1
      rom[1138] = 8'b00111100;  // 2   ****
      rom[1139] = 8'b01100110;  // 3  **  **
      rom[1140] = 8'b11000010;  // 4 **    *
      rom[1141] = 8'b11000000;  // 5 **
      rom[1142] = 8'b11000000;  // 6 **
      rom[1143] = 8'b11011110;  // 7 ** ****
      rom[1144] = 8'b11000110;  // 8 **   **
      rom[1145] = 8'b11000110;  // 9 **   **
      rom[1146] = 8'b01100110;  // a  **  **
      rom[1147] = 8'b00111010;  // b   *** *
      rom[1148] = 8'b00000000;  // c
      rom[1149] = 8'b00000000;  // d
      rom[1150] = 8'b00000000;  // e
      rom[1151] = 8'b00000000;  // f
      // code x48
      rom[1152] = 8'b00000000;  // 0
      rom[1153] = 8'b00000000;  // 1
      rom[1154] = 8'b11000110;  // 2 **   **
      rom[1155] = 8'b11000110;  // 3 **   **
      rom[1156] = 8'b11000110;  // 4 **   **
      rom[1157] = 8'b11000110;  // 5 **   **
      rom[1158] = 8'b11111110;  // 6 *******
      rom[1159] = 8'b11000110;  // 7 **   **
      rom[1160] = 8'b11000110;  // 8 **   **
      rom[1161] = 8'b11000110;  // 9 **   **
      rom[1162] = 8'b11000110;  // a **   **
      rom[1163] = 8'b11000110;  // b **   **
      rom[1164] = 8'b00000000;  // c
      rom[1165] = 8'b00000000;  // d
      rom[1166] = 8'b00000000;  // e
      rom[1167] = 8'b00000000;  // f
      // code x49
      rom[1168] = 8'b00000000;  // 0
      rom[1169] = 8'b00000000;  // 1
      rom[1170] = 8'b00111100;  // 2   ****
      rom[1171] = 8'b00011000;  // 3    **
      rom[1172] = 8'b00011000;  // 4    **
      rom[1173] = 8'b00011000;  // 5    **
      rom[1174] = 8'b00011000;  // 6    **
      rom[1175] = 8'b00011000;  // 7    **
      rom[1176] = 8'b00011000;  // 8    **
      rom[1177] = 8'b00011000;  // 9    **
      rom[1178] = 8'b00011000;  // a    **
      rom[1179] = 8'b00111100;  // b   ****
      rom[1180] = 8'b00000000;  // c
      rom[1181] = 8'b00000000;  // d
      rom[1182] = 8'b00000000;  // e
      rom[1183] = 8'b00000000;  // f
      // code x4a
      rom[1184] = 8'b00000000;  // 0
      rom[1185] = 8'b00000000;  // 1
      rom[1186] = 8'b00011110;  // 2    ****
      rom[1187] = 8'b00001100;  // 3     **
      rom[1188] = 8'b00001100;  // 4     **
      rom[1189] = 8'b00001100;  // 5     **
      rom[1190] = 8'b00001100;  // 6     **
      rom[1191] = 8'b00001100;  // 7     **
      rom[1192] = 8'b11001100;  // 8 **  **
      rom[1193] = 8'b11001100;  // 9 **  **
      rom[1194] = 8'b11001100;  // a **  **
      rom[1195] = 8'b01111000;  // b  ****
      rom[1196] = 8'b00000000;  // c
      rom[1197] = 8'b00000000;  // d
      rom[1198] = 8'b00000000;  // e
      rom[1199] = 8'b00000000;  // f
      // code x4b
      rom[1200] = 8'b00000000;  // 0
      rom[1201] = 8'b00000000;  // 1
      rom[1202] = 8'b11100110;  // 2 ***  **
      rom[1203] = 8'b01100110;  // 3  **  **
      rom[1204] = 8'b01100110;  // 4  **  **
      rom[1205] = 8'b01101100;  // 5  ** **
      rom[1206] = 8'b01111000;  // 6  ****
      rom[1207] = 8'b01111000;  // 7  ****
      rom[1208] = 8'b01101100;  // 8  ** **
      rom[1209] = 8'b01100110;  // 9  **  **
      rom[1210] = 8'b01100110;  // a  **  **
      rom[1211] = 8'b11100110;  // b ***  **
      rom[1212] = 8'b00000000;  // c
      rom[1213] = 8'b00000000;  // d
      rom[1214] = 8'b00000000;  // e
      rom[1215] = 8'b00000000;  // f
      // code x4c
      rom[1216] = 8'b00000000;  // 0
      rom[1217] = 8'b00000000;  // 1
      rom[1218] = 8'b11110000;  // 2 ****
      rom[1219] = 8'b01100000;  // 3  **
      rom[1220] = 8'b01100000;  // 4  **
      rom[1221] = 8'b01100000;  // 5  **
      rom[1222] = 8'b01100000;  // 6  **
      rom[1223] = 8'b01100000;  // 7  **
      rom[1224] = 8'b01100000;  // 8  **
      rom[1225] = 8'b01100010;  // 9  **   *
      rom[1226] = 8'b01100110;  // a  **  **
      rom[1227] = 8'b11111110;  // b *******
      rom[1228] = 8'b00000000;  // c
      rom[1229] = 8'b00000000;  // d
      rom[1230] = 8'b00000000;  // e
      rom[1231] = 8'b00000000;  // f
      // code x4d
      rom[1232] = 8'b00000000;  // 0
      rom[1233] = 8'b00000000;  // 1
      rom[1234] = 8'b11000011;  // 2 **    **
      rom[1235] = 8'b11100111;  // 3 ***  ***
      rom[1236] = 8'b11111111;  // 4 ********
      rom[1237] = 8'b11111111;  // 5 ********
      rom[1238] = 8'b11011011;  // 6 ** ** **
      rom[1239] = 8'b11000011;  // 7 **    **
      rom[1240] = 8'b11000011;  // 8 **    **
      rom[1241] = 8'b11000011;  // 9 **    **
      rom[1242] = 8'b11000011;  // a **    **
      rom[1243] = 8'b11000011;  // b **    **
      rom[1244] = 8'b00000000;  // c
      rom[1245] = 8'b00000000;  // d
      rom[1246] = 8'b00000000;  // e
      rom[1247] = 8'b00000000;  // f
      // code x4e
      rom[1248] = 8'b00000000;  // 0
      rom[1249] = 8'b00000000;  // 1
      rom[1250] = 8'b11000110;  // 2 **   **
      rom[1251] = 8'b11100110;  // 3 ***  **
      rom[1252] = 8'b11110110;  // 4 **** **
      rom[1253] = 8'b11111110;  // 5 *******
      rom[1254] = 8'b11011110;  // 6 ** ****
      rom[1255] = 8'b11001110;  // 7 **  ***
      rom[1256] = 8'b11000110;  // 8 **   **
      rom[1257] = 8'b11000110;  // 9 **   **
      rom[1258] = 8'b11000110;  // a **   **
      rom[1259] = 8'b11000110;  // b **   **
      rom[1260] = 8'b00000000;  // c
      rom[1261] = 8'b00000000;  // d
      rom[1262] = 8'b00000000;  // e
      rom[1263] = 8'b00000000;  // f
      // code x4f
      rom[1264] = 8'b00000000;  // 0
      rom[1265] = 8'b00000000;  // 1
      rom[1266] = 8'b01111100;  // 2  *****
      rom[1267] = 8'b11000110;  // 3 **   **
      rom[1268] = 8'b11000110;  // 4 **   **
      rom[1269] = 8'b11000110;  // 5 **   **
      rom[1270] = 8'b11000110;  // 6 **   **
      rom[1271] = 8'b11000110;  // 7 **   **
      rom[1272] = 8'b11000110;  // 8 **   **
      rom[1273] = 8'b11000110;  // 9 **   **
      rom[1274] = 8'b11000110;  // a **   **
      rom[1275] = 8'b01111100;  // b  *****
      rom[1276] = 8'b00000000;  // c
      rom[1277] = 8'b00000000;  // d
      rom[1278] = 8'b00000000;  // e
      rom[1279] = 8'b00000000;  // f
      // code x50
      rom[1280] = 8'b00000000;  // 0
      rom[1281] = 8'b00000000;  // 1
      rom[1282] = 8'b11111100;  // 2 ******
      rom[1283] = 8'b01100110;  // 3  **  **
      rom[1284] = 8'b01100110;  // 4  **  **
      rom[1285] = 8'b01100110;  // 5  **  **
      rom[1286] = 8'b01111100;  // 6  *****
      rom[1287] = 8'b01100000;  // 7  **
      rom[1288] = 8'b01100000;  // 8  **
      rom[1289] = 8'b01100000;  // 9  **
      rom[1290] = 8'b01100000;  // a  **
      rom[1291] = 8'b11110000;  // b ****
      rom[1292] = 8'b00000000;  // c
      rom[1293] = 8'b00000000;  // d
      rom[1294] = 8'b00000000;  // e
      rom[1295] = 8'b00000000;  // f
      // code x510
      rom[1296] = 8'b00000000;  // 0
      rom[1297] = 8'b00000000;  // 1
      rom[1298] = 8'b01111100;  // 2  *****
      rom[1299] = 8'b11000110;  // 3 **   **
      rom[1300] = 8'b11000110;  // 4 **   **
      rom[1301] = 8'b11000110;  // 5 **   **
      rom[1302] = 8'b11000110;  // 6 **   **
      rom[1303] = 8'b11000110;  // 7 **   **
      rom[1304] = 8'b11000110;  // 8 **   **
      rom[1305] = 8'b11010110;  // 9 ** * **
      rom[1306] = 8'b11011110;  // a ** ****
      rom[1307] = 8'b01111100;  // b  *****
      rom[1308] = 8'b00001100;  // c     **
      rom[1309] = 8'b00001110;  // d     ***
      rom[1310] = 8'b00000000;  // e
      rom[1311] = 8'b00000000;  // f
      // code x52
      rom[1312] = 8'b00000000;  // 0
      rom[1313] = 8'b00000000;  // 1
      rom[1314] = 8'b11111100;  // 2 ******
      rom[1315] = 8'b01100110;  // 3  **  **
      rom[1316] = 8'b01100110;  // 4  **  **
      rom[1317] = 8'b01100110;  // 5  **  **
      rom[1318] = 8'b01111100;  // 6  *****
      rom[1319] = 8'b01101100;  // 7  ** **
      rom[1320] = 8'b01100110;  // 8  **  **
      rom[1321] = 8'b01100110;  // 9  **  **
      rom[1322] = 8'b01100110;  // a  **  **
      rom[1323] = 8'b11100110;  // b ***  **
      rom[1324] = 8'b00000000;  // c
      rom[1325] = 8'b00000000;  // d
      rom[1326] = 8'b00000000;  // e
      rom[1327] = 8'b00000000;  // f
      // code x53
      rom[1328] = 8'b00000000;  // 0
      rom[1329] = 8'b00000000;  // 1
      rom[1330] = 8'b01111100;  // 2  *****
      rom[1331] = 8'b11000110;  // 3 **   **
      rom[1332] = 8'b11000110;  // 4 **   **
      rom[1333] = 8'b01100000;  // 5  **
      rom[1334] = 8'b00111000;  // 6   ***
      rom[1335] = 8'b00001100;  // 7     **
      rom[1336] = 8'b00000110;  // 8      **
      rom[1337] = 8'b11000110;  // 9 **   **
      rom[1338] = 8'b11000110;  // a **   **
      rom[1339] = 8'b01111100;  // b  *****
      rom[1340] = 8'b00000000;  // c
      rom[1341] = 8'b00000000;  // d
      rom[1342] = 8'b00000000;  // e
      rom[1343] = 8'b00000000;  // f
      // code x54
      rom[1344] = 8'b00000000;  // 0
      rom[1345] = 8'b00000000;  // 1
      rom[1346] = 8'b11111111;  // 2 ********
      rom[1347] = 8'b11011011;  // 3 ** ** **
      rom[1348] = 8'b10011001;  // 4 *  **  *
      rom[1349] = 8'b00011000;  // 5    **
      rom[1350] = 8'b00011000;  // 6    **
      rom[1351] = 8'b00011000;  // 7    **
      rom[1352] = 8'b00011000;  // 8    **
      rom[1353] = 8'b00011000;  // 9    **
      rom[1354] = 8'b00011000;  // a    **
      rom[1355] = 8'b00111100;  // b   ****
      rom[1356] = 8'b00000000;  // c
      rom[1357] = 8'b00000000;  // d
      rom[1358] = 8'b00000000;  // e
      rom[1359] = 8'b00000000;  // f
      // code x55
      rom[1360] = 8'b00000000;  // 0
      rom[1361] = 8'b00000000;  // 1
      rom[1362] = 8'b11000110;  // 2 **   **
      rom[1363] = 8'b11000110;  // 3 **   **
      rom[1364] = 8'b11000110;  // 4 **   **
      rom[1365] = 8'b11000110;  // 5 **   **
      rom[1366] = 8'b11000110;  // 6 **   **
      rom[1367] = 8'b11000110;  // 7 **   **
      rom[1368] = 8'b11000110;  // 8 **   **
      rom[1369] = 8'b11000110;  // 9 **   **
      rom[1370] = 8'b11000110;  // a **   **
      rom[1371] = 8'b01111100;  // b  *****
      rom[1372] = 8'b00000000;  // c
      rom[1373] = 8'b00000000;  // d
      rom[1374] = 8'b00000000;  // e
      rom[1375] = 8'b00000000;  // f
      // code x56
      rom[1376] = 8'b00000000;  // 0
      rom[1377] = 8'b00000000;  // 1
      rom[1378] = 8'b11000011;  // 2 **    **
      rom[1379] = 8'b11000011;  // 3 **    **
      rom[1380] = 8'b11000011;  // 4 **    **
      rom[1381] = 8'b11000011;  // 5 **    **
      rom[1382] = 8'b11000011;  // 6 **    **
      rom[1383] = 8'b11000011;  // 7 **    **
      rom[1384] = 8'b11000011;  // 8 **    **
      rom[1385] = 8'b01100110;  // 9  **  **
      rom[1386] = 8'b00111100;  // a   ****
      rom[1387] = 8'b00011000;  // b    **
      rom[1388] = 8'b00000000;  // c
      rom[1389] = 8'b00000000;  // d
      rom[1390] = 8'b00000000;  // e
      rom[1391] = 8'b00000000;  // f
      // code x57
      rom[1392] = 8'b00000000;  // 0
      rom[1393] = 8'b00000000;  // 1
      rom[1394] = 8'b11000011;  // 2 **    **
      rom[1395] = 8'b11000011;  // 3 **    **
      rom[1396] = 8'b11000011;  // 4 **    **
      rom[1397] = 8'b11000011;  // 5 **    **
      rom[1398] = 8'b11000011;  // 6 **    **
      rom[1399] = 8'b11011011;  // 7 ** ** **
      rom[1400] = 8'b11011011;  // 8 ** ** **
      rom[1401] = 8'b11111111;  // 9 ********
      rom[1402] = 8'b01100110;  // a  **  **
      rom[1403] = 8'b01100110;  // b  **  **
      rom[1404] = 8'b00000000;  // c
      rom[1405] = 8'b00000000;  // d
      rom[1406] = 8'b00000000;  // e
      rom[1407] = 8'b00000000;  // f

      // code x58
      rom[1408] = 8'b00000000;  // 0
      rom[1409] = 8'b00000000;  // 1
      rom[1410] = 8'b11000011;  // 2 **    **
      rom[1411] = 8'b11000011;  // 3 **    **
      rom[1412] = 8'b01100110;  // 4  **  **
      rom[1413] = 8'b00111100;  // 5   ****
      rom[1414] = 8'b00011000;  // 6    **
      rom[1415] = 8'b00011000;  // 7    **
      rom[1416] = 8'b00111100;  // 8   ****
      rom[1417] = 8'b01100110;  // 9  **  **
      rom[1418] = 8'b11000011;  // a **    **
      rom[1419] = 8'b11000011;  // b **    **
      rom[1420] = 8'b00000000;  // c
      rom[1421] = 8'b00000000;  // d
      rom[1422] = 8'b00000000;  // e
      rom[1423] = 8'b00000000;  // f
      // code x59
      rom[1424] = 8'b00000000;  // 0
      rom[1425] = 8'b00000000;  // 1
      rom[1426] = 8'b11000011;  // 2 **    **
      rom[1427] = 8'b11000011;  // 3 **    **
      rom[1428] = 8'b11000011;  // 4 **    **
      rom[1429] = 8'b01100110;  // 5  **  **
      rom[1430] = 8'b00111100;  // 6   ****
      rom[1431] = 8'b00011000;  // 7    **
      rom[1432] = 8'b00011000;  // 8    **
      rom[1433] = 8'b00011000;  // 9    **
      rom[1434] = 8'b00011000;  // a    **
      rom[1435] = 8'b00111100;  // b   ****
      rom[1436] = 8'b00000000;  // c
      rom[1437] = 8'b00000000;  // d
      rom[1438] = 8'b00000000;  // e
      rom[1439] = 8'b00000000;  // f
      // code x5a
      rom[1440] = 8'b00000000;  // 0
      rom[1441] = 8'b00000000;  // 1
      rom[1442] = 8'b11111111;  // 2 ********
      rom[1443] = 8'b11000011;  // 3 **    **
      rom[1444] = 8'b10000110;  // 4 *    **
      rom[1445] = 8'b00001100;  // 5     **
      rom[1446] = 8'b00011000;  // 6    **
      rom[1447] = 8'b00110000;  // 7   **
      rom[1448] = 8'b01100000;  // 8  **
      rom[1449] = 8'b11000001;  // 9 **     *
      rom[1450] = 8'b11000011;  // a **    **
      rom[1451] = 8'b11111111;  // b ********
      rom[1452] = 8'b00000000;  // c
      rom[1453] = 8'b00000000;  // d
      rom[1454] = 8'b00000000;  // e
      rom[1455] = 8'b00000000;  // f
      // code x5b
      rom[1456] = 8'b00000000;  // 0
      rom[1457] = 8'b00000000;  // 1
      rom[1458] = 8'b00111100;  // 2   ****
      rom[1459] = 8'b00110000;  // 3   **
      rom[1460] = 8'b00110000;  // 4   **
      rom[1461] = 8'b00110000;  // 5   **
      rom[1462] = 8'b00110000;  // 6   **
      rom[1463] = 8'b00110000;  // 7   **
      rom[1464] = 8'b00110000;  // 8   **
      rom[1465] = 8'b00110000;  // 9   **
      rom[1466] = 8'b00110000;  // a   **
      rom[1467] = 8'b00111100;  // b   ****
      rom[1468] = 8'b00000000;  // c
      rom[1469] = 8'b00000000;  // d
      rom[1470] = 8'b00000000;  // e
      rom[1471] = 8'b00000000;  // f
      // code x5c
      rom[1472] = 8'b00000000;  // 0
      rom[1473] = 8'b00000000;  // 1
      rom[1474] = 8'b00000000;  // 2
      rom[1475] = 8'b10000000;  // 3 *
      rom[1476] = 8'b11000000;  // 4 **
      rom[1477] = 8'b11100000;  // 5 ***
      rom[1478] = 8'b01110000;  // 6  ***
      rom[1479] = 8'b00111000;  // 7   ***
      rom[1480] = 8'b00011100;  // 8    ***
      rom[1481] = 8'b00001110;  // 9     ***
      rom[1482] = 8'b00000110;  // a      **
      rom[1483] = 8'b00000010;  // b       *
      rom[1484] = 8'b00000000;  // c
      rom[1485] = 8'b00000000;  // d
      rom[1486] = 8'b00000000;  // e
      rom[1487] = 8'b00000000;  // f
      // code x5d
      rom[1488] = 8'b00000000;  // 0
      rom[1489] = 8'b00000000;  // 1
      rom[1490] = 8'b00111100;  // 2   ****
      rom[1491] = 8'b00001100;  // 3     **
      rom[1492] = 8'b00001100;  // 4     **
      rom[1493] = 8'b00001100;  // 5     **
      rom[1494] = 8'b00001100;  // 6     **
      rom[1495] = 8'b00001100;  // 7     **
      rom[1496] = 8'b00001100;  // 8     **
      rom[1497] = 8'b00001100;  // 9     **
      rom[1498] = 8'b00001100;  // a     **
      rom[1499] = 8'b00111100;  // b   ****
      rom[1500] = 8'b00000000;  // c
      rom[1501] = 8'b00000000;  // d
      rom[1502] = 8'b00000000;  // e
      rom[1503] = 8'b00000000;  // f
      // code x5e
      rom[1504] = 8'b00010000;  // 0    *
      rom[1505] = 8'b00111000;  // 1   ***
      rom[1506] = 8'b01101100;  // 2  ** **
      rom[1507] = 8'b11000110;  // 3 **   **
      rom[1508] = 8'b00000000;  // 4
      rom[1509] = 8'b00000000;  // 5
      rom[1510] = 8'b00000000;  // 6
      rom[1511] = 8'b00000000;  // 7
      rom[1512] = 8'b00000000;  // 8
      rom[1513] = 8'b00000000;  // 9
      rom[1514] = 8'b00000000;  // a
      rom[1515] = 8'b00000000;  // b
      rom[1516] = 8'b00000000;  // c
      rom[1517] = 8'b00000000;  // d
      rom[1518] = 8'b00000000;  // e
      rom[1519] = 8'b00000000;  // f
      // code x5f
      rom[1520] = 8'b00000000;  // 0
      rom[1521] = 8'b00000000;  // 1
      rom[1522] = 8'b00000000;  // 2
      rom[1523] = 8'b00000000;  // 3
      rom[1524] = 8'b00000000;  // 4
      rom[1525] = 8'b00000000;  // 5
      rom[1526] = 8'b00000000;  // 6
      rom[1527] = 8'b00000000;  // 7
      rom[1528] = 8'b00000000;  // 8
      rom[1529] = 8'b00000000;  // 9
      rom[1530] = 8'b00000000;  // a
      rom[1531] = 8'b00000000;  // b
      rom[1532] = 8'b00000000;  // c
      rom[1533] = 8'b11111111;  // d ********
      rom[1534] = 8'b00000000;  // e
      rom[1535] = 8'b00000000;  // f
      // code x60
      rom[1536] = 8'b00110000;  // 0   **
      rom[1537] = 8'b00110000;  // 1   **
      rom[1538] = 8'b00011000;  // 2    **
      rom[1539] = 8'b00000000;  // 3
      rom[1540] = 8'b00000000;  // 4
      rom[1541] = 8'b00000000;  // 5
      rom[1542] = 8'b00000000;  // 6
      rom[1543] = 8'b00000000;  // 7
      rom[1544] = 8'b00000000;  // 8
      rom[1545] = 8'b00000000;  // 9
      rom[1546] = 8'b00000000;  // a
      rom[1547] = 8'b00000000;  // b
      rom[1548] = 8'b00000000;  // c
      rom[1549] = 8'b00000000;  // d
      rom[1550] = 8'b00000000;  // e
      rom[1551] = 8'b00000000;  // f
      // code x61
      rom[1552] = 8'b00000000;  // 0
      rom[1553] = 8'b00000000;  // 1
      rom[1554] = 8'b00000000;  // 2
      rom[1555] = 8'b00000000;  // 3
      rom[1556] = 8'b00000000;  // 4
      rom[1557] = 8'b01111000;  // 5  ****
      rom[1558] = 8'b00001100;  // 6     **
      rom[1559] = 8'b01111100;  // 7  *****
      rom[1560] = 8'b11001100;  // 8 **  **
      rom[1561] = 8'b11001100;  // 9 **  **
      rom[1562] = 8'b11001100;  // a **  **
      rom[1563] = 8'b01110110;  // b  *** **
      rom[1564] = 8'b00000000;  // c
      rom[1565] = 8'b00000000;  // d
      rom[1566] = 8'b00000000;  // e
      rom[1567] = 8'b00000000;  // f
      // code x62
      rom[1568] = 8'b00000000;  // 0
      rom[1569] = 8'b00000000;  // 1
      rom[1570] = 8'b11100000;  // 2  ***
      rom[1571] = 8'b01100000;  // 3   **
      rom[1572] = 8'b01100000;  // 4   **
      rom[1573] = 8'b01111000;  // 5   ****
      rom[1574] = 8'b01101100;  // 6   ** **
      rom[1575] = 8'b01100110;  // 7   **  **
      rom[1576] = 8'b01100110;  // 8   **  **
      rom[1577] = 8'b01100110;  // 9   **  **
      rom[1578] = 8'b01100110;  // a   **  **
      rom[1579] = 8'b01111100;  // b   *****
      rom[1580] = 8'b00000000;  // c
      rom[1581] = 8'b00000000;  // d
      rom[1582] = 8'b00000000;  // e
      rom[1583] = 8'b00000000;  // f
      // code x63
      rom[1584] = 8'b00000000;  // 0
      rom[1585] = 8'b00000000;  // 1
      rom[1586] = 8'b00000000;  // 2
      rom[1587] = 8'b00000000;  // 3
      rom[1588] = 8'b00000000;  // 4
      rom[1589] = 8'b01111100;  // 5  *****
      rom[1590] = 8'b11000110;  // 6 **   **
      rom[1591] = 8'b11000000;  // 7 **
      rom[1592] = 8'b11000000;  // 8 **
      rom[1593] = 8'b11000000;  // 9 **
      rom[1594] = 8'b11000110;  // a **   **
      rom[1595] = 8'b01111100;  // b  *****
      rom[1596] = 8'b00000000;  // c
      rom[1597] = 8'b00000000;  // d
      rom[1598] = 8'b00000000;  // e
      rom[1599] = 8'b00000000;  // f
      // code x64
      rom[1600] = 8'b00000000;  // 0
      rom[1601] = 8'b00000000;  // 1
      rom[1602] = 8'b00011100;  // 2    ***
      rom[1603] = 8'b00001100;  // 3     **
      rom[1604] = 8'b00001100;  // 4     **
      rom[1605] = 8'b00111100;  // 5   ****
      rom[1606] = 8'b01101100;  // 6  ** **
      rom[1607] = 8'b11001100;  // 7 **  **
      rom[1608] = 8'b11001100;  // 8 **  **
      rom[1609] = 8'b11001100;  // 9 **  **
      rom[1610] = 8'b11001100;  // a **  **
      rom[1611] = 8'b01110110;  // b  *** **
      rom[1612] = 8'b00000000;  // c
      rom[1613] = 8'b00000000;  // d
      rom[1614] = 8'b00000000;  // e
      rom[1615] = 8'b00000000;  // f
      // code x65
      rom[1616] = 8'b00000000;  // 0
      rom[1617] = 8'b00000000;  // 1
      rom[1618] = 8'b00000000;  // 2
      rom[1619] = 8'b00000000;  // 3
      rom[1620] = 8'b00000000;  // 4
      rom[1621] = 8'b01111100;  // 5  *****
      rom[1622] = 8'b11000110;  // 6 **   **
      rom[1623] = 8'b11111110;  // 7 *******
      rom[1624] = 8'b11000000;  // 8 **
      rom[1625] = 8'b11000000;  // 9 **
      rom[1626] = 8'b11000110;  // a **   **
      rom[1627] = 8'b01111100;  // b  *****
      rom[1628] = 8'b00000000;  // c
      rom[1629] = 8'b00000000;  // d
      rom[1630] = 8'b00000000;  // e
      rom[1631] = 8'b00000000;  // f
      // code x66
      rom[1632] = 8'b00000000;  // 0
      rom[1633] = 8'b00000000;  // 1
      rom[1634] = 8'b00111000;  // 2   ***
      rom[1635] = 8'b01101100;  // 3  ** **
      rom[1636] = 8'b01100100;  // 4  **  *
      rom[1637] = 8'b01100000;  // 5  **
      rom[1638] = 8'b11110000;  // 6 ****
      rom[1639] = 8'b01100000;  // 7  **
      rom[1640] = 8'b01100000;  // 8  **
      rom[1641] = 8'b01100000;  // 9  **
      rom[1642] = 8'b01100000;  // a  **
      rom[1643] = 8'b11110000;  // b ****
      rom[1644] = 8'b00000000;  // c
      rom[1645] = 8'b00000000;  // d
      rom[1646] = 8'b00000000;  // e
      rom[1647] = 8'b00000000;  // f
      // code x67
      rom[1648] = 8'b00000000;  // 0
      rom[1649] = 8'b00000000;  // 1
      rom[1650] = 8'b00000000;  // 2
      rom[1651] = 8'b00000000;  // 3
      rom[1652] = 8'b00000000;  // 4
      rom[1653] = 8'b01110110;  // 5  *** **
      rom[1654] = 8'b11001100;  // 6 **  **
      rom[1655] = 8'b11001100;  // 7 **  **
      rom[1656] = 8'b11001100;  // 8 **  **
      rom[1657] = 8'b11001100;  // 9 **  **
      rom[1658] = 8'b11001100;  // a **  **
      rom[1659] = 8'b01111100;  // b  *****
      rom[1660] = 8'b00001100;  // c     **
      rom[1661] = 8'b11001100;  // d **  **
      rom[1662] = 8'b01111000;  // e  ****
      rom[1663] = 8'b00000000;  // f
      // code x68
      rom[1664] = 8'b00000000;  // 0
      rom[1665] = 8'b00000000;  // 1
      rom[1666] = 8'b11100000;  // 2 ***
      rom[1667] = 8'b01100000;  // 3  **
      rom[1668] = 8'b01100000;  // 4  **
      rom[1669] = 8'b01101100;  // 5  ** **
      rom[1670] = 8'b01110110;  // 6  *** **
      rom[1671] = 8'b01100110;  // 7  **  **
      rom[1672] = 8'b01100110;  // 8  **  **
      rom[1673] = 8'b01100110;  // 9  **  **
      rom[1674] = 8'b01100110;  // a  **  **
      rom[1675] = 8'b11100110;  // b ***  **
      rom[1676] = 8'b00000000;  // c
      rom[1677] = 8'b00000000;  // d
      rom[1678] = 8'b00000000;  // e
      rom[1679] = 8'b00000000;  // f
      // code x69
      rom[1680] = 8'b00000000;  // 0
      rom[1681] = 8'b00000000;  // 1
      rom[1682] = 8'b00011000;  // 2    **
      rom[1683] = 8'b00011000;  // 3    **
      rom[1684] = 8'b00000000;  // 4
      rom[1685] = 8'b00111000;  // 5   ***
      rom[1686] = 8'b00011000;  // 6    **
      rom[1687] = 8'b00011000;  // 7    **
      rom[1688] = 8'b00011000;  // 8    **
      rom[1689] = 8'b00011000;  // 9    **
      rom[1690] = 8'b00011000;  // a    **
      rom[1691] = 8'b00111100;  // b   ****
      rom[1692] = 8'b00000000;  // c
      rom[1693] = 8'b00000000;  // d
      rom[1694] = 8'b00000000;  // e
      rom[1695] = 8'b00000000;  // f
      // code x6a
      rom[1696] = 8'b00000000;  // 0
      rom[1697] = 8'b00000000;  // 1
      rom[1698] = 8'b00000110;  // 2      **
      rom[1699] = 8'b00000110;  // 3      **
      rom[1700] = 8'b00000000;  // 4
      rom[1701] = 8'b00001110;  // 5     ***
      rom[1702] = 8'b00000110;  // 6      **
      rom[1703] = 8'b00000110;  // 7      **
      rom[1704] = 8'b00000110;  // 8      **
      rom[1705] = 8'b00000110;  // 9      **
      rom[1706] = 8'b00000110;  // a      **
      rom[1707] = 8'b00000110;  // b      **
      rom[1708] = 8'b01100110;  // c  **  **
      rom[1709] = 8'b01100110;  // d  **  **
      rom[1710] = 8'b00111100;  // e   ****
      rom[1711] = 8'b00000000;  // f
      // code x6b
      rom[1712] = 8'b00000000;  // 0
      rom[1713] = 8'b00000000;  // 1
      rom[1714] = 8'b11100000;  // 2 ***
      rom[1715] = 8'b01100000;  // 3  **
      rom[1716] = 8'b01100000;  // 4  **
      rom[1717] = 8'b01100110;  // 5  **  **
      rom[1718] = 8'b01101100;  // 6  ** **
      rom[1719] = 8'b01111000;  // 7  ****
      rom[1720] = 8'b01111000;  // 8  ****
      rom[1721] = 8'b01101100;  // 9  ** **
      rom[1722] = 8'b01100110;  // a  **  **
      rom[1723] = 8'b11100110;  // b ***  **
      rom[1724] = 8'b00000000;  // c
      rom[1725] = 8'b00000000;  // d
      rom[1726] = 8'b00000000;  // e
      rom[1727] = 8'b00000000;  // f
      // code x6c
      rom[1728] = 8'b00000000;  // 0
      rom[1729] = 8'b00000000;  // 1
      rom[1730] = 8'b00111000;  // 2   ***
      rom[1731] = 8'b00011000;  // 3    **
      rom[1732] = 8'b00011000;  // 4    **
      rom[1733] = 8'b00011000;  // 5    **
      rom[1734] = 8'b00011000;  // 6    **
      rom[1735] = 8'b00011000;  // 7    **
      rom[1736] = 8'b00011000;  // 8    **
      rom[1737] = 8'b00011000;  // 9    **
      rom[1738] = 8'b00011000;  // a    **
      rom[1739] = 8'b00111100;  // b   ****
      rom[1740] = 8'b00000000;  // c
      rom[1741] = 8'b00000000;  // d
      rom[1742] = 8'b00000000;  // e
      rom[1743] = 8'b00000000;  // f
      // code x6d
      rom[1744] = 8'b00000000;  // 0
      rom[1745] = 8'b00000000;  // 1
      rom[1746] = 8'b00000000;  // 2
      rom[1747] = 8'b00000000;  // 3
      rom[1748] = 8'b00000000;  // 4
      rom[1749] = 8'b11100110;  // 5 ***  **
      rom[1750] = 8'b11111111;  // 6 ********
      rom[1751] = 8'b11011011;  // 7 ** ** **
      rom[1752] = 8'b11011011;  // 8 ** ** **
      rom[1753] = 8'b11011011;  // 9 ** ** **
      rom[1754] = 8'b11011011;  // a ** ** **
      rom[1755] = 8'b11011011;  // b ** ** **
      rom[1756] = 8'b00000000;  // c
      rom[1757] = 8'b00000000;  // d
      rom[1758] = 8'b00000000;  // e
      rom[1759] = 8'b00000000;  // f
      // code x6e
      rom[1760] = 8'b00000000;  // 0
      rom[1761] = 8'b00000000;  // 1
      rom[1762] = 8'b00000000;  // 2
      rom[1763] = 8'b00000000;  // 3
      rom[1764] = 8'b00000000;  // 4
      rom[1765] = 8'b11011100;  // 5 ** ***
      rom[1766] = 8'b01100110;  // 6  **  **
      rom[1767] = 8'b01100110;  // 7  **  **
      rom[1768] = 8'b01100110;  // 8  **  **
      rom[1769] = 8'b01100110;  // 9  **  **
      rom[1770] = 8'b01100110;  // a  **  **
      rom[1771] = 8'b01100110;  // b  **  **
      rom[1772] = 8'b00000000;  // c
      rom[1773] = 8'b00000000;  // d
      rom[1774] = 8'b00000000;  // e
      rom[1775] = 8'b00000000;  // f
      // code x6f
      rom[1776] = 8'b00000000;  // 0
      rom[1777] = 8'b00000000;  // 1
      rom[1778] = 8'b00000000;  // 2
      rom[1779] = 8'b00000000;  // 3
      rom[1780] = 8'b00000000;  // 4
      rom[1781] = 8'b01111100;  // 5  *****
      rom[1782] = 8'b11000110;  // 6 **   **
      rom[1783] = 8'b11000110;  // 7 **   **
      rom[1784] = 8'b11000110;  // 8 **   **
      rom[1785] = 8'b11000110;  // 9 **   **
      rom[1786] = 8'b11000110;  // a **   **
      rom[1787] = 8'b01111100;  // b  *****
      rom[1788] = 8'b00000000;  // c
      rom[1789] = 8'b00000000;  // d
      rom[1790] = 8'b00000000;  // e
      rom[1791] = 8'b00000000;  // f
      // code x70
      rom[1792] = 8'b00000000;  // 0
      rom[1793] = 8'b00000000;  // 1
      rom[1794] = 8'b00000000;  // 2
      rom[1795] = 8'b00000000;  // 3
      rom[1796] = 8'b00000000;  // 4
      rom[1797] = 8'b11011100;  // 5 ** ***
      rom[1798] = 8'b01100110;  // 6  **  **
      rom[1799] = 8'b01100110;  // 7  **  **
      rom[1800] = 8'b01100110;  // 8  **  **
      rom[1801] = 8'b01100110;  // 9  **  **
      rom[1802] = 8'b01100110;  // a  **  **
      rom[1803] = 8'b01111100;  // b  *****
      rom[1804] = 8'b01100000;  // c  **
      rom[1805] = 8'b01100000;  // d  **
      rom[1806] = 8'b11110000;  // e ****
      rom[1807] = 8'b00000000;  // f
      // code x71
      rom[1808] = 8'b00000000;  // 0
      rom[1809] = 8'b00000000;  // 1
      rom[1810] = 8'b00000000;  // 2
      rom[1811] = 8'b00000000;  // 3
      rom[1812] = 8'b00000000;  // 4
      rom[1813] = 8'b01110110;  // 5  *** **
      rom[1814] = 8'b11001100;  // 6 **  **
      rom[1815] = 8'b11001100;  // 7 **  **
      rom[1816] = 8'b11001100;  // 8 **  **
      rom[1817] = 8'b11001100;  // 9 **  **
      rom[1818] = 8'b11001100;  // a **  **
      rom[1819] = 8'b01111100;  // b  *****
      rom[1820] = 8'b00001100;  // c     **
      rom[1821] = 8'b00001100;  // d     **
      rom[1822] = 8'b00011110;  // e    ****
      rom[1823] = 8'b00000000;  // f
      // code x72
      rom[1824] = 8'b00000000;  // 0
      rom[1825] = 8'b00000000;  // 1
      rom[1826] = 8'b00000000;  // 2
      rom[1827] = 8'b00000000;  // 3
      rom[1828] = 8'b00000000;  // 4
      rom[1829] = 8'b11011100;  // 5 ** ***
      rom[1830] = 8'b01110110;  // 6  *** **
      rom[1831] = 8'b01100110;  // 7  **  **
      rom[1832] = 8'b01100000;  // 8  **
      rom[1833] = 8'b01100000;  // 9  **
      rom[1834] = 8'b01100000;  // a  **
      rom[1835] = 8'b11110000;  // b ****
      rom[1836] = 8'b00000000;  // c
      rom[1837] = 8'b00000000;  // d
      rom[1838] = 8'b00000000;  // e
      rom[1839] = 8'b00000000;  // f
      // code x73
      rom[1840] = 8'b00000000;  // 0
      rom[1841] = 8'b00000000;  // 1
      rom[1842] = 8'b00000000;  // 2
      rom[1843] = 8'b00000000;  // 3
      rom[1844] = 8'b00000000;  // 4
      rom[1845] = 8'b01111100;  // 5  *****
      rom[1846] = 8'b11000110;  // 6 **   **
      rom[1847] = 8'b01100000;  // 7  **
      rom[1848] = 8'b00111000;  // 8   ***
      rom[1849] = 8'b00001100;  // 9     **
      rom[1850] = 8'b11000110;  // a **   **
      rom[1851] = 8'b01111100;  // b  *****
      rom[1852] = 8'b00000000;  // c
      rom[1853] = 8'b00000000;  // d
      rom[1854] = 8'b00000000;  // e
      rom[1855] = 8'b00000000;  // f
      // code x74
      rom[1856] = 8'b00000000;  // 0
      rom[1857] = 8'b00000000;  // 1
      rom[1858] = 8'b00010000;  // 2    *
      rom[1859] = 8'b00110000;  // 3   **
      rom[1860] = 8'b00110000;  // 4   **
      rom[1861] = 8'b11111100;  // 5 ******
      rom[1862] = 8'b00110000;  // 6   **
      rom[1863] = 8'b00110000;  // 7   **
      rom[1864] = 8'b00110000;  // 8   **
      rom[1865] = 8'b00110000;  // 9   **
      rom[1866] = 8'b00110110;  // a   ** **
      rom[1867] = 8'b00011100;  // b    ***
      rom[1868] = 8'b00000000;  // c
      rom[1869] = 8'b00000000;  // d
      rom[1870] = 8'b00000000;  // e
      rom[1871] = 8'b00000000;  // f
      // code x75
      rom[1872] = 8'b00000000;  // 0
      rom[1873] = 8'b00000000;  // 1
      rom[1874] = 8'b00000000;  // 2
      rom[1875] = 8'b00000000;  // 3
      rom[1876] = 8'b00000000;  // 4
      rom[1877] = 8'b11001100;  // 5 **  **
      rom[1878] = 8'b11001100;  // 6 **  **
      rom[1879] = 8'b11001100;  // 7 **  **
      rom[1880] = 8'b11001100;  // 8 **  **
      rom[1881] = 8'b11001100;  // 9 **  **
      rom[1882] = 8'b11001100;  // a **  **
      rom[1883] = 8'b01110110;  // b  *** **
      rom[1884] = 8'b00000000;  // c
      rom[1885] = 8'b00000000;  // d
      rom[1886] = 8'b00000000;  // e
      rom[1887] = 8'b00000000;  // f
      // code x76
      rom[1888] = 8'b00000000;  // 0
      rom[1889] = 8'b00000000;  // 1
      rom[1890] = 8'b00000000;  // 2
      rom[1891] = 8'b00000000;  // 3
      rom[1892] = 8'b00000000;  // 4
      rom[1893] = 8'b11000011;  // 5 **    **
      rom[1894] = 8'b11000011;  // 6 **    **
      rom[1895] = 8'b11000011;  // 7 **    **
      rom[1896] = 8'b11000011;  // 8 **    **
      rom[1897] = 8'b01100110;  // 9  **  **
      rom[1898] = 8'b00111100;  // a   ****
      rom[1899] = 8'b00011000;  // b    **
      rom[1900] = 8'b00000000;  // c
      rom[1901] = 8'b00000000;  // d
      rom[1902] = 8'b00000000;  // e
      rom[1903] = 8'b00000000;  // f
      // code x77
      rom[1904] = 8'b00000000;  // 0
      rom[1905] = 8'b00000000;  // 1
      rom[1906] = 8'b00000000;  // 2
      rom[1907] = 8'b00000000;  // 3
      rom[1908] = 8'b00000000;  // 4
      rom[1909] = 8'b11000011;  // 5 **    **
      rom[1910] = 8'b11000011;  // 6 **    **
      rom[1911] = 8'b11000011;  // 7 **    **
      rom[1912] = 8'b11011011;  // 8 ** ** **
      rom[1913] = 8'b11011011;  // 9 ** ** **
      rom[1914] = 8'b11111111;  // a ********
      rom[1915] = 8'b01100110;  // b  **  **
      rom[1916] = 8'b00000000;  // c
      rom[1917] = 8'b00000000;  // d
      rom[1918] = 8'b00000000;  // e
      rom[1919] = 8'b00000000;  // f
      // code x78
      rom[1920] = 8'b00000000;  // 0
      rom[1921] = 8'b00000000;  // 1
      rom[1922] = 8'b00000000;  // 2
      rom[1923] = 8'b00000000;  // 3
      rom[1924] = 8'b00000000;  // 4
      rom[1925] = 8'b11000011;  // 5 **    **
      rom[1926] = 8'b01100110;  // 6  **  **
      rom[1927] = 8'b00111100;  // 7   ****
      rom[1928] = 8'b00011000;  // 8    **
      rom[1929] = 8'b00111100;  // 9   ****
      rom[1930] = 8'b01100110;  // a  **  **
      rom[1931] = 8'b11000011;  // b **    **
      rom[1932] = 8'b00000000;  // c
      rom[1933] = 8'b00000000;  // d
      rom[1934] = 8'b00000000;  // e
      rom[1935] = 8'b00000000;  // f
      // code x79
      rom[1936] = 8'b00000000;  // 0
      rom[1937] = 8'b00000000;  // 1
      rom[1938] = 8'b00000000;  // 2
      rom[1939] = 8'b00000000;  // 3
      rom[1940] = 8'b00000000;  // 4
      rom[1941] = 8'b11000110;  // 5 **   **
      rom[1942] = 8'b11000110;  // 6 **   **
      rom[1943] = 8'b11000110;  // 7 **   **
      rom[1944] = 8'b11000110;  // 8 **   **
      rom[1945] = 8'b11000110;  // 9 **   **
      rom[1946] = 8'b11000110;  // a **   **
      rom[1947] = 8'b01111110;  // b  ******
      rom[1948] = 8'b00000110;  // c      **
      rom[1949] = 8'b00001100;  // d     **
      rom[1950] = 8'b11111000;  // e *****
      rom[1951] = 8'b00000000;  // f
      // code x7a
      rom[1952] = 8'b00000000;  // 0
      rom[1953] = 8'b00000000;  // 1
      rom[1954] = 8'b00000000;  // 2
      rom[1955] = 8'b00000000;  // 3
      rom[1956] = 8'b00000000;  // 4
      rom[1957] = 8'b11111110;  // 5 *******
      rom[1958] = 8'b11001100;  // 6 **  **
      rom[1959] = 8'b00011000;  // 7    **
      rom[1960] = 8'b00110000;  // 8   **
      rom[1961] = 8'b01100000;  // 9  **
      rom[1962] = 8'b11000110;  // a **   **
      rom[1963] = 8'b11111110;  // b *******
      rom[1964] = 8'b00000000;  // c
      rom[1965] = 8'b00000000;  // d
      rom[1966] = 8'b00000000;  // e
      rom[1967] = 8'b00000000;  // f
      // code x7b
      rom[1968] = 8'b00000000;  // 0
      rom[1969] = 8'b00000000;  // 1
      rom[1970] = 8'b00001110;  // 2     ***
      rom[1971] = 8'b00011000;  // 3    **
      rom[1972] = 8'b00011000;  // 4    **
      rom[1973] = 8'b00011000;  // 5    **
      rom[1974] = 8'b01110000;  // 6  ***
      rom[1975] = 8'b00011000;  // 7    **
      rom[1976] = 8'b00011000;  // 8    **
      rom[1977] = 8'b00011000;  // 9    **
      rom[1978] = 8'b00011000;  // a    **
      rom[1979] = 8'b00001110;  // b     ***
      rom[1980] = 8'b00000000;  // c
      rom[1981] = 8'b00000000;  // d
      rom[1982] = 8'b00000000;  // e
      rom[1983] = 8'b00000000;  // f
      // code x7c
      rom[1984] = 8'b00000000;  // 0
      rom[1985] = 8'b00000000;  // 1
      rom[1986] = 8'b00011000;  // 2    **
      rom[1987] = 8'b00011000;  // 3    **
      rom[1988] = 8'b00011000;  // 4    **
      rom[1989] = 8'b00011000;  // 5    **
      rom[1990] = 8'b00000000;  // 6
      rom[1991] = 8'b00011000;  // 7    **
      rom[1992] = 8'b00011000;  // 8    **
      rom[1993] = 8'b00011000;  // 9    **
      rom[1994] = 8'b00011000;  // a    **
      rom[1995] = 8'b00011000;  // b    **
      rom[1996] = 8'b00000000;  // c
      rom[1997] = 8'b00000000;  // d
      rom[1998] = 8'b00000000;  // e
      rom[1999] = 8'b00000000;  // f
      // code x7d
      rom[2000] = 8'b00000000;  // 0
      rom[2001] = 8'b00000000;  // 1
      rom[2002] = 8'b01110000;  // 2  ***
      rom[2003] = 8'b00011000;  // 3    **
      rom[2004] = 8'b00011000;  // 4    **
      rom[2005] = 8'b00011000;  // 5    **
      rom[2006] = 8'b00001110;  // 6     ***
      rom[2007] = 8'b00011000;  // 7    **
      rom[2008] = 8'b00011000;  // 8    **
      rom[2009] = 8'b00011000;  // 9    **
      rom[2010] = 8'b00011000;  // a    **
      rom[2011] = 8'b01110000;  // b  ***
      rom[2012] = 8'b00000000;  // c
      rom[2013] = 8'b00000000;  // d
      rom[2014] = 8'b00000000;  // e
      rom[2015] = 8'b00000000;  // f
      // code x7e
      rom[2016] = 8'b00000000;  // 0
      rom[2017] = 8'b00000000;  // 1
      rom[2018] = 8'b01110110;  // 2  *** **
      rom[2019] = 8'b11011100;  // 3 ** ***
      rom[2020] = 8'b00000000;  // 4
      rom[2021] = 8'b00000000;  // 5
      rom[2022] = 8'b00000000;  // 6
      rom[2023] = 8'b00000000;  // 7
      rom[2024] = 8'b00000000;  // 8
      rom[2025] = 8'b00000000;  // 9
      rom[2026] = 8'b00000000;  // a
      rom[2027] = 8'b00000000;  // b
      rom[2028] = 8'b00000000;  // c
      rom[2029] = 8'b00000000;  // d
      rom[2030] = 8'b00000000;  // e
      rom[2031] = 8'b00000000;  // f
      // code x7f
      rom[2032] = 8'b00000000;  // 0
      rom[2033] = 8'b00000000;  // 1
      rom[2034] = 8'b00000000;  // 2
      rom[2035] = 8'b00000000;  // 3
      rom[2036] = 8'b00010000;  // 4    *
      rom[2037] = 8'b00111000;  // 5   ***
      rom[2038] = 8'b01101100;  // 6  ** **
      rom[2039] = 8'b11000110;  // 7 **   **
      rom[2040] = 8'b11000110;  // 8 **   **
      rom[2041] = 8'b11000110;  // 9 **   **
      rom[2042] = 8'b11111110;  // a *******
      rom[2043] = 8'b00000000;  // b
      rom[2044] = 8'b00000000;  // c
      rom[2045] = 8'b00000000;  // d
      rom[2046] = 8'b00000000;  // e
      rom[2047] = 8'b00000000;  // f
   end

   always_ff @(posedge clk)
      addr_reg <= addr;

   assign data = rom[addr_reg];

endmodule



